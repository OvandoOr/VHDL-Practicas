library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM_Chirp is
   port(
      CLK : in std_logic;
      I   : in  std_logic_vector(9 downto 0);
      A   : out std_logic_vector(7 downto 0)
      );
   end entity;

architecture ROM of ROM_Chirp is

subtype word_t is std_logic_vector(7 downto 0);
type memory_t is array(0 to 1023) of word_t;

signal rom : memory_t := (         -- Coefficient format 1.7
   "00100010", -- Column 1   Coefficient 0.26562500
   "00100011", -- Column 2   Coefficient 0.27343750
   "00100010", -- Column 3   Coefficient 0.26562500
   "00100010", -- Column 4   Coefficient 0.26562500
   "00100001", -- Column 5   Coefficient 0.25781250
   "00100001", -- Column 6   Coefficient 0.25781250
   "00100001", -- Column 7   Coefficient 0.25781250
   "00100010", -- Column 8   Coefficient 0.26562500
   "00100010", -- Column 9   Coefficient 0.26562500
   "00100001", -- Column 10   Coefficient 0.25781250
   "00100001", -- Column 11   Coefficient 0.25781250
   "00100001", -- Column 12   Coefficient 0.25781250
   "00100001", -- Column 13   Coefficient 0.25781250
   "00100001", -- Column 14   Coefficient 0.25781250
   "00100000", -- Column 15   Coefficient 0.25000000
   "00100000", -- Column 16   Coefficient 0.25000000
   "00100001", -- Column 17   Coefficient 0.25781250
   "00100001", -- Column 18   Coefficient 0.25781250
   "00100001", -- Column 19   Coefficient 0.25781250
   "00100001", -- Column 20   Coefficient 0.25781250
   "00100000", -- Column 21   Coefficient 0.25000000
   "00100001", -- Column 22   Coefficient 0.25781250
   "00100001", -- Column 23   Coefficient 0.25781250
   "00100001", -- Column 24   Coefficient 0.25781250
   "00100001", -- Column 25   Coefficient 0.25781250
   "00100001", -- Column 26   Coefficient 0.25781250
   "00100000", -- Column 27   Coefficient 0.25000000
   "00100000", -- Column 28   Coefficient 0.25000000
   "00100001", -- Column 29   Coefficient 0.25781250
   "00100001", -- Column 30   Coefficient 0.25781250
   "00100001", -- Column 31   Coefficient 0.25781250
   "00100000", -- Column 32   Coefficient 0.25000000
   "00100000", -- Column 33   Coefficient 0.25000000
   "00100001", -- Column 34   Coefficient 0.25781250
   "00100001", -- Column 35   Coefficient 0.25781250
   "00100001", -- Column 36   Coefficient 0.25781250
   "00100001", -- Column 37   Coefficient 0.25781250
   "00100001", -- Column 38   Coefficient 0.25781250
   "00100001", -- Column 39   Coefficient 0.25781250
   "00100000", -- Column 40   Coefficient 0.25000000
   "00100000", -- Column 41   Coefficient 0.25000000
   "00100000", -- Column 42   Coefficient 0.25000000
   "00100000", -- Column 43   Coefficient 0.25000000
   "00100000", -- Column 44   Coefficient 0.25000000
   "00100000", -- Column 45   Coefficient 0.25000000
   "00011111", -- Column 46   Coefficient 0.24218750
   "00011111", -- Column 47   Coefficient 0.24218750
   "00100000", -- Column 48   Coefficient 0.25000000
   "00100000", -- Column 49   Coefficient 0.25000000
   "00100000", -- Column 50   Coefficient 0.25000000
   "00011111", -- Column 51   Coefficient 0.24218750
   "00011111", -- Column 52   Coefficient 0.24218750
   "00011111", -- Column 53   Coefficient 0.24218750
   "00100000", -- Column 54   Coefficient 0.25000000
   "00100000", -- Column 55   Coefficient 0.25000000
   "00100000", -- Column 56   Coefficient 0.25000000
   "00100000", -- Column 57   Coefficient 0.25000000
   "00100000", -- Column 58   Coefficient 0.25000000
   "00011111", -- Column 59   Coefficient 0.24218750
   "00011111", -- Column 60   Coefficient 0.24218750
   "00011111", -- Column 61   Coefficient 0.24218750
   "00100000", -- Column 62   Coefficient 0.25000000
   "00100000", -- Column 63   Coefficient 0.25000000
   "00100000", -- Column 64   Coefficient 0.25000000
   "00100000", -- Column 65   Coefficient 0.25000000
   "00100000", -- Column 66   Coefficient 0.25000000
   "00011111", -- Column 67   Coefficient 0.24218750
   "00100000", -- Column 68   Coefficient 0.25000000
   "00100000", -- Column 69   Coefficient 0.25000000
   "00100000", -- Column 70   Coefficient 0.25000000
   "00100000", -- Column 71   Coefficient 0.25000000
   "00100000", -- Column 72   Coefficient 0.25000000
   "00100000", -- Column 73   Coefficient 0.25000000
   "00100000", -- Column 74   Coefficient 0.25000000
   "00100000", -- Column 75   Coefficient 0.25000000
   "00100000", -- Column 76   Coefficient 0.25000000
   "00100000", -- Column 77   Coefficient 0.25000000
   "00100000", -- Column 78   Coefficient 0.25000000
   "00100001", -- Column 79   Coefficient 0.25781250
   "00100000", -- Column 80   Coefficient 0.25000000
   "00100000", -- Column 81   Coefficient 0.25000000
   "00100000", -- Column 82   Coefficient 0.25000000
   "00100000", -- Column 83   Coefficient 0.25000000
   "00100000", -- Column 84   Coefficient 0.25000000
   "00100001", -- Column 85   Coefficient 0.25781250
   "00100010", -- Column 86   Coefficient 0.26562500
   "00100010", -- Column 87   Coefficient 0.26562500
   "00100010", -- Column 88   Coefficient 0.26562500
   "00100010", -- Column 89   Coefficient 0.26562500
   "00100010", -- Column 90   Coefficient 0.26562500
   "00100010", -- Column 91   Coefficient 0.26562500
   "00100001", -- Column 92   Coefficient 0.25781250
   "00100010", -- Column 93   Coefficient 0.26562500
   "00100011", -- Column 94   Coefficient 0.27343750
   "00100011", -- Column 95   Coefficient 0.27343750
   "00100011", -- Column 96   Coefficient 0.27343750
   "00100011", -- Column 97   Coefficient 0.27343750
   "00100100", -- Column 98   Coefficient 0.28125000
   "00100101", -- Column 99   Coefficient 0.28906250
   "00100110", -- Column 100   Coefficient 0.29687500
   "00100110", -- Column 101   Coefficient 0.29687500
   "00100110", -- Column 102   Coefficient 0.29687500
   "00100110", -- Column 103   Coefficient 0.29687500
   "00100110", -- Column 104   Coefficient 0.29687500
   "00100110", -- Column 105   Coefficient 0.29687500
   "00100111", -- Column 106   Coefficient 0.30468750
   "00100111", -- Column 107   Coefficient 0.30468750
   "00100111", -- Column 108   Coefficient 0.30468750
   "00101000", -- Column 109   Coefficient 0.31250000
   "00101000", -- Column 110   Coefficient 0.31250000
   "00101000", -- Column 111   Coefficient 0.31250000
   "00101000", -- Column 112   Coefficient 0.31250000
   "00101000", -- Column 113   Coefficient 0.31250000
   "00101000", -- Column 114   Coefficient 0.31250000
   "00101000", -- Column 115   Coefficient 0.31250000
   "00101000", -- Column 116   Coefficient 0.31250000
   "00101000", -- Column 117   Coefficient 0.31250000
   "00101001", -- Column 118   Coefficient 0.32031250
   "00101001", -- Column 119   Coefficient 0.32031250
   "00101010", -- Column 120   Coefficient 0.32812500
   "00101010", -- Column 121   Coefficient 0.32812500
   "00101010", -- Column 122   Coefficient 0.32812500
   "00101011", -- Column 123   Coefficient 0.33593750
   "00101011", -- Column 124   Coefficient 0.33593750
   "00101011", -- Column 125   Coefficient 0.33593750
   "00101011", -- Column 126   Coefficient 0.33593750
   "00101011", -- Column 127   Coefficient 0.33593750
   "00101011", -- Column 128   Coefficient 0.33593750
   "00101100", -- Column 129   Coefficient 0.34375000
   "00101100", -- Column 130   Coefficient 0.34375000
   "00101100", -- Column 131   Coefficient 0.34375000
   "00101011", -- Column 132   Coefficient 0.33593750
   "00101011", -- Column 133   Coefficient 0.33593750
   "00101100", -- Column 134   Coefficient 0.34375000
   "00101100", -- Column 135   Coefficient 0.34375000
   "00101100", -- Column 136   Coefficient 0.34375000
   "00101100", -- Column 137   Coefficient 0.34375000
   "00101011", -- Column 138   Coefficient 0.33593750
   "00101011", -- Column 139   Coefficient 0.33593750
   "00101011", -- Column 140   Coefficient 0.33593750
   "00101011", -- Column 141   Coefficient 0.33593750
   "00101011", -- Column 142   Coefficient 0.33593750
   "00101011", -- Column 143   Coefficient 0.33593750
   "00101011", -- Column 144   Coefficient 0.33593750
   "00101011", -- Column 145   Coefficient 0.33593750
   "00101011", -- Column 146   Coefficient 0.33593750
   "00101011", -- Column 147   Coefficient 0.33593750
   "00101100", -- Column 148   Coefficient 0.34375000
   "00101100", -- Column 149   Coefficient 0.34375000
   "00101100", -- Column 150   Coefficient 0.34375000
   "00101100", -- Column 151   Coefficient 0.34375000
   "00101100", -- Column 152   Coefficient 0.34375000
   "00101011", -- Column 153   Coefficient 0.33593750
   "00101010", -- Column 154   Coefficient 0.32812500
   "00101001", -- Column 155   Coefficient 0.32031250
   "00101001", -- Column 156   Coefficient 0.32031250
   "00101010", -- Column 157   Coefficient 0.32812500
   "00101010", -- Column 158   Coefficient 0.32812500
   "00101010", -- Column 159   Coefficient 0.32812500
   "00101011", -- Column 160   Coefficient 0.33593750
   "00101011", -- Column 161   Coefficient 0.33593750
   "00101011", -- Column 162   Coefficient 0.33593750
   "00101010", -- Column 163   Coefficient 0.32812500
   "00101010", -- Column 164   Coefficient 0.32812500
   "00101010", -- Column 165   Coefficient 0.32812500
   "00101010", -- Column 166   Coefficient 0.32812500
   "00101001", -- Column 167   Coefficient 0.32031250
   "00101001", -- Column 168   Coefficient 0.32031250
   "00101000", -- Column 169   Coefficient 0.31250000
   "00100111", -- Column 170   Coefficient 0.30468750
   "00100110", -- Column 171   Coefficient 0.29687500
   "00100100", -- Column 172   Coefficient 0.28125000
   "00100100", -- Column 173   Coefficient 0.28125000
   "00100011", -- Column 174   Coefficient 0.27343750
   "00100011", -- Column 175   Coefficient 0.27343750
   "00100010", -- Column 176   Coefficient 0.26562500
   "00100001", -- Column 177   Coefficient 0.25781250
   "00100001", -- Column 178   Coefficient 0.25781250
   "00100001", -- Column 179   Coefficient 0.25781250
   "00100001", -- Column 180   Coefficient 0.25781250
   "00100000", -- Column 181   Coefficient 0.25000000
   "00011111", -- Column 182   Coefficient 0.24218750
   "00011111", -- Column 183   Coefficient 0.24218750
   "00011111", -- Column 184   Coefficient 0.24218750
   "00011111", -- Column 185   Coefficient 0.24218750
   "00011110", -- Column 186   Coefficient 0.23437500
   "00011111", -- Column 187   Coefficient 0.24218750
   "00100000", -- Column 188   Coefficient 0.25000000
   "00100000", -- Column 189   Coefficient 0.25000000
   "00100000", -- Column 190   Coefficient 0.25000000
   "00100000", -- Column 191   Coefficient 0.25000000
   "00100000", -- Column 192   Coefficient 0.25000000
   "00100000", -- Column 193   Coefficient 0.25000000
   "00011111", -- Column 194   Coefficient 0.24218750
   "00011111", -- Column 195   Coefficient 0.24218750
   "00011111", -- Column 196   Coefficient 0.24218750
   "00100000", -- Column 197   Coefficient 0.25000000
   "00100000", -- Column 198   Coefficient 0.25000000
   "00011111", -- Column 199   Coefficient 0.24218750
   "00011110", -- Column 200   Coefficient 0.23437500
   "00011111", -- Column 201   Coefficient 0.24218750
   "00011110", -- Column 202   Coefficient 0.23437500
   "00011101", -- Column 203   Coefficient 0.22656250
   "00011100", -- Column 204   Coefficient 0.21875000
   "00011101", -- Column 205   Coefficient 0.22656250
   "00011101", -- Column 206   Coefficient 0.22656250
   "00011101", -- Column 207   Coefficient 0.22656250
   "00011101", -- Column 208   Coefficient 0.22656250
   "00011110", -- Column 209   Coefficient 0.23437500
   "00011110", -- Column 210   Coefficient 0.23437500
   "00011110", -- Column 211   Coefficient 0.23437500
   "00011101", -- Column 212   Coefficient 0.22656250
   "00011100", -- Column 213   Coefficient 0.21875000
   "00011101", -- Column 214   Coefficient 0.22656250
   "00011101", -- Column 215   Coefficient 0.22656250
   "00011101", -- Column 216   Coefficient 0.22656250
   "00011101", -- Column 217   Coefficient 0.22656250
   "00011101", -- Column 218   Coefficient 0.22656250
   "00011101", -- Column 219   Coefficient 0.22656250
   "00011100", -- Column 220   Coefficient 0.21875000
   "00011100", -- Column 221   Coefficient 0.21875000
   "00011100", -- Column 222   Coefficient 0.21875000
   "00011101", -- Column 223   Coefficient 0.22656250
   "00011101", -- Column 224   Coefficient 0.22656250
   "00011101", -- Column 225   Coefficient 0.22656250
   "00011101", -- Column 226   Coefficient 0.22656250
   "00011101", -- Column 227   Coefficient 0.22656250
   "00011101", -- Column 228   Coefficient 0.22656250
   "00011101", -- Column 229   Coefficient 0.22656250
   "00011100", -- Column 230   Coefficient 0.21875000
   "00011101", -- Column 231   Coefficient 0.22656250
   "00011101", -- Column 232   Coefficient 0.22656250
   "00011110", -- Column 233   Coefficient 0.23437500
   "00011110", -- Column 234   Coefficient 0.23437500
   "00011101", -- Column 235   Coefficient 0.22656250
   "00011101", -- Column 236   Coefficient 0.22656250
   "00011101", -- Column 237   Coefficient 0.22656250
   "00011110", -- Column 238   Coefficient 0.23437500
   "00011110", -- Column 239   Coefficient 0.23437500
   "00011110", -- Column 240   Coefficient 0.23437500
   "00011110", -- Column 241   Coefficient 0.23437500
   "00011110", -- Column 242   Coefficient 0.23437500
   "00011110", -- Column 243   Coefficient 0.23437500
   "00011101", -- Column 244   Coefficient 0.22656250
   "00011101", -- Column 245   Coefficient 0.22656250
   "00011101", -- Column 246   Coefficient 0.22656250
   "00011110", -- Column 247   Coefficient 0.23437500
   "00011111", -- Column 248   Coefficient 0.24218750
   "00011110", -- Column 249   Coefficient 0.23437500
   "00011110", -- Column 250   Coefficient 0.23437500
   "00011110", -- Column 251   Coefficient 0.23437500
   "00011110", -- Column 252   Coefficient 0.23437500
   "00011110", -- Column 253   Coefficient 0.23437500
   "00011110", -- Column 254   Coefficient 0.23437500
   "00011110", -- Column 255   Coefficient 0.23437500
   "00011111", -- Column 256   Coefficient 0.24218750
   "00011110", -- Column 257   Coefficient 0.23437500
   "00011101", -- Column 258   Coefficient 0.22656250
   "00011101", -- Column 259   Coefficient 0.22656250
   "00011110", -- Column 260   Coefficient 0.23437500
   "00011110", -- Column 261   Coefficient 0.23437500
   "00011110", -- Column 262   Coefficient 0.23437500
   "00011111", -- Column 263   Coefficient 0.24218750
   "00100001", -- Column 264   Coefficient 0.25781250
   "00100010", -- Column 265   Coefficient 0.26562500
   "00100011", -- Column 266   Coefficient 0.27343750
   "00100100", -- Column 267   Coefficient 0.28125000
   "00100111", -- Column 268   Coefficient 0.30468750
   "00101001", -- Column 269   Coefficient 0.32031250
   "00101100", -- Column 270   Coefficient 0.34375000
   "00101111", -- Column 271   Coefficient 0.36718750
   "00110010", -- Column 272   Coefficient 0.39062500
   "00110101", -- Column 273   Coefficient 0.41406250
   "00111000", -- Column 274   Coefficient 0.43750000
   "00111100", -- Column 275   Coefficient 0.46875000
   "01000011", -- Column 276   Coefficient 0.52343750
   "01001011", -- Column 277   Coefficient 0.58593750
   "01010010", -- Column 278   Coefficient 0.64062500
   "01011010", -- Column 279   Coefficient 0.70312500
   "01100010", -- Column 280   Coefficient 0.76562500
   "01101010", -- Column 281   Coefficient 0.82812500
   "01110010", -- Column 282   Coefficient 0.89062500
   "01111001", -- Column 283   Coefficient 0.94531250
   "01111100", -- Column 284   Coefficient 0.96875000
   "01111101", -- Column 285   Coefficient 0.97656250
   "01111101", -- Column 286   Coefficient 0.97656250
   "01111100", -- Column 287   Coefficient 0.96875000
   "01111101", -- Column 288   Coefficient 0.97656250
   "01111111", -- Column 289   Coefficient 0.99218750
   "01111110", -- Column 290   Coefficient 0.98437500
   "01111011", -- Column 291   Coefficient 0.96093750
   "01111000", -- Column 292   Coefficient 0.93750000
   "01110111", -- Column 293   Coefficient 0.92968750
   "01110111", -- Column 294   Coefficient 0.92968750
   "01110110", -- Column 295   Coefficient 0.92187500
   "01110011", -- Column 296   Coefficient 0.89843750
   "01110000", -- Column 297   Coefficient 0.87500000
   "01101110", -- Column 298   Coefficient 0.85937500
   "01101011", -- Column 299   Coefficient 0.83593750
   "01100111", -- Column 300   Coefficient 0.80468750
   "01100011", -- Column 301   Coefficient 0.77343750
   "01100001", -- Column 302   Coefficient 0.75781250
   "01011110", -- Column 303   Coefficient 0.73437500
   "01010111", -- Column 304   Coefficient 0.67968750
   "01001110", -- Column 305   Coefficient 0.60937500
   "01000111", -- Column 306   Coefficient 0.55468750
   "01000011", -- Column 307   Coefficient 0.52343750
   "00111110", -- Column 308   Coefficient 0.48437500
   "00110001", -- Column 309   Coefficient 0.38281250
   "00011101", -- Column 310   Coefficient 0.22656250
   "00001011", -- Column 311   Coefficient 0.08593750
   "00000100", -- Column 312   Coefficient 0.03125000
   "00000101", -- Column 313   Coefficient 0.03906250
   "00000111", -- Column 314   Coefficient 0.05468750
   "00000111", -- Column 315   Coefficient 0.05468750
   "00001000", -- Column 316   Coefficient 0.06250000
   "00001100", -- Column 317   Coefficient 0.09375000
   "00001111", -- Column 318   Coefficient 0.11718750
   "00010001", -- Column 319   Coefficient 0.13281250
   "00010011", -- Column 320   Coefficient 0.14843750
   "00010110", -- Column 321   Coefficient 0.17187500
   "00011010", -- Column 322   Coefficient 0.20312500
   "00011110", -- Column 323   Coefficient 0.23437500
   "00100010", -- Column 324   Coefficient 0.26562500
   "00100101", -- Column 325   Coefficient 0.28906250
   "00101000", -- Column 326   Coefficient 0.31250000
   "00101001", -- Column 327   Coefficient 0.32031250
   "00101010", -- Column 328   Coefficient 0.32812500
   "00101011", -- Column 329   Coefficient 0.33593750
   "00101011", -- Column 330   Coefficient 0.33593750
   "00101101", -- Column 331   Coefficient 0.35156250
   "00101110", -- Column 332   Coefficient 0.35937500
   "00110000", -- Column 333   Coefficient 0.37500000
   "00110001", -- Column 334   Coefficient 0.38281250
   "00110001", -- Column 335   Coefficient 0.38281250
   "00110001", -- Column 336   Coefficient 0.38281250
   "00110010", -- Column 337   Coefficient 0.39062500
   "00110010", -- Column 338   Coefficient 0.39062500
   "00110011", -- Column 339   Coefficient 0.39843750
   "00110011", -- Column 340   Coefficient 0.39843750
   "00110011", -- Column 341   Coefficient 0.39843750
   "00110011", -- Column 342   Coefficient 0.39843750
   "00110011", -- Column 343   Coefficient 0.39843750
   "00110011", -- Column 344   Coefficient 0.39843750
   "00110100", -- Column 345   Coefficient 0.40625000
   "00110100", -- Column 346   Coefficient 0.40625000
   "00110011", -- Column 347   Coefficient 0.39843750
   "00110011", -- Column 348   Coefficient 0.39843750
   "00110100", -- Column 349   Coefficient 0.40625000
   "00110100", -- Column 350   Coefficient 0.40625000
   "00110100", -- Column 351   Coefficient 0.40625000
   "00110011", -- Column 352   Coefficient 0.39843750
   "00110011", -- Column 353   Coefficient 0.39843750
   "00110011", -- Column 354   Coefficient 0.39843750
   "00110011", -- Column 355   Coefficient 0.39843750
   "00110011", -- Column 356   Coefficient 0.39843750
   "00110011", -- Column 357   Coefficient 0.39843750
   "00110011", -- Column 358   Coefficient 0.39843750
   "00110011", -- Column 359   Coefficient 0.39843750
   "00110100", -- Column 360   Coefficient 0.40625000
   "00110101", -- Column 361   Coefficient 0.41406250
   "00110101", -- Column 362   Coefficient 0.41406250
   "00110101", -- Column 363   Coefficient 0.41406250
   "00110101", -- Column 364   Coefficient 0.41406250
   "00110101", -- Column 365   Coefficient 0.41406250
   "00110101", -- Column 366   Coefficient 0.41406250
   "00110101", -- Column 367   Coefficient 0.41406250
   "00110101", -- Column 368   Coefficient 0.41406250
   "00110110", -- Column 369   Coefficient 0.42187500
   "00110110", -- Column 370   Coefficient 0.42187500
   "00110111", -- Column 371   Coefficient 0.42968750
   "00110110", -- Column 372   Coefficient 0.42187500
   "00110110", -- Column 373   Coefficient 0.42187500
   "00110111", -- Column 374   Coefficient 0.42968750
   "00110111", -- Column 375   Coefficient 0.42968750
   "00110111", -- Column 376   Coefficient 0.42968750
   "00111000", -- Column 377   Coefficient 0.43750000
   "00111000", -- Column 378   Coefficient 0.43750000
   "00111000", -- Column 379   Coefficient 0.43750000
   "00110111", -- Column 380   Coefficient 0.42968750
   "00110111", -- Column 381   Coefficient 0.42968750
   "00111000", -- Column 382   Coefficient 0.43750000
   "00111000", -- Column 383   Coefficient 0.43750000
   "00110111", -- Column 384   Coefficient 0.42968750
   "00111000", -- Column 385   Coefficient 0.43750000
   "00111001", -- Column 386   Coefficient 0.44531250
   "00111010", -- Column 387   Coefficient 0.45312500
   "00111010", -- Column 388   Coefficient 0.45312500
   "00111010", -- Column 389   Coefficient 0.45312500
   "00111010", -- Column 390   Coefficient 0.45312500
   "00111010", -- Column 391   Coefficient 0.45312500
   "00111010", -- Column 392   Coefficient 0.45312500
   "00111010", -- Column 393   Coefficient 0.45312500
   "00111011", -- Column 394   Coefficient 0.46093750
   "00111100", -- Column 395   Coefficient 0.46875000
   "00111100", -- Column 396   Coefficient 0.46875000
   "00111011", -- Column 397   Coefficient 0.46093750
   "00111011", -- Column 398   Coefficient 0.46093750
   "00111100", -- Column 399   Coefficient 0.46875000
   "00111100", -- Column 400   Coefficient 0.46875000
   "00111100", -- Column 401   Coefficient 0.46875000
   "00111100", -- Column 402   Coefficient 0.46875000
   "00111101", -- Column 403   Coefficient 0.47656250
   "00111101", -- Column 404   Coefficient 0.47656250
   "00111100", -- Column 405   Coefficient 0.46875000
   "00111100", -- Column 406   Coefficient 0.46875000
   "00111101", -- Column 407   Coefficient 0.47656250
   "00111110", -- Column 408   Coefficient 0.48437500
   "00111110", -- Column 409   Coefficient 0.48437500
   "00111110", -- Column 410   Coefficient 0.48437500
   "00111110", -- Column 411   Coefficient 0.48437500
   "00111110", -- Column 412   Coefficient 0.48437500
   "00111110", -- Column 413   Coefficient 0.48437500
   "00111110", -- Column 414   Coefficient 0.48437500
   "00111110", -- Column 415   Coefficient 0.48437500
   "00111110", -- Column 416   Coefficient 0.48437500
   "00111111", -- Column 417   Coefficient 0.49218750
   "00111111", -- Column 418   Coefficient 0.49218750
   "01000000", -- Column 419   Coefficient 0.50000000
   "01000000", -- Column 420   Coefficient 0.50000000
   "01000001", -- Column 421   Coefficient 0.50781250
   "01000000", -- Column 422   Coefficient 0.50000000
   "01000001", -- Column 423   Coefficient 0.50781250
   "01000000", -- Column 424   Coefficient 0.50000000
   "01000001", -- Column 425   Coefficient 0.50781250
   "01000001", -- Column 426   Coefficient 0.50781250
   "01000001", -- Column 427   Coefficient 0.50781250
   "01000010", -- Column 428   Coefficient 0.51562500
   "01000010", -- Column 429   Coefficient 0.51562500
   "01000011", -- Column 430   Coefficient 0.52343750
   "01000011", -- Column 431   Coefficient 0.52343750
   "01000010", -- Column 432   Coefficient 0.51562500
   "01000010", -- Column 433   Coefficient 0.51562500
   "01000011", -- Column 434   Coefficient 0.52343750
   "01000100", -- Column 435   Coefficient 0.53125000
   "01000101", -- Column 436   Coefficient 0.53906250
   "01000101", -- Column 437   Coefficient 0.53906250
   "01000101", -- Column 438   Coefficient 0.53906250
   "01000110", -- Column 439   Coefficient 0.54687500
   "01000101", -- Column 440   Coefficient 0.53906250
   "01000110", -- Column 441   Coefficient 0.54687500
   "01000110", -- Column 442   Coefficient 0.54687500
   "01000110", -- Column 443   Coefficient 0.54687500
   "01000110", -- Column 444   Coefficient 0.54687500
   "01000110", -- Column 445   Coefficient 0.54687500
   "01000111", -- Column 446   Coefficient 0.55468750
   "01001000", -- Column 447   Coefficient 0.56250000
   "01001000", -- Column 448   Coefficient 0.56250000
   "01001000", -- Column 449   Coefficient 0.56250000
   "01000111", -- Column 450   Coefficient 0.55468750
   "01001000", -- Column 451   Coefficient 0.56250000
   "01001000", -- Column 452   Coefficient 0.56250000
   "01001000", -- Column 453   Coefficient 0.56250000
   "01001001", -- Column 454   Coefficient 0.57031250
   "01001001", -- Column 455   Coefficient 0.57031250
   "01001001", -- Column 456   Coefficient 0.57031250
   "01001001", -- Column 457   Coefficient 0.57031250
   "01001001", -- Column 458   Coefficient 0.57031250
   "01001010", -- Column 459   Coefficient 0.57812500
   "01001011", -- Column 460   Coefficient 0.58593750
   "01001011", -- Column 461   Coefficient 0.58593750
   "01001011", -- Column 462   Coefficient 0.58593750
   "01001011", -- Column 463   Coefficient 0.58593750
   "01001100", -- Column 464   Coefficient 0.59375000
   "01001100", -- Column 465   Coefficient 0.59375000
   "01001100", -- Column 466   Coefficient 0.59375000
   "01001101", -- Column 467   Coefficient 0.60156250
   "01001101", -- Column 468   Coefficient 0.60156250
   "01001101", -- Column 469   Coefficient 0.60156250
   "01001101", -- Column 470   Coefficient 0.60156250
   "01001111", -- Column 471   Coefficient 0.61718750
   "01001111", -- Column 472   Coefficient 0.61718750
   "01001111", -- Column 473   Coefficient 0.61718750
   "01001110", -- Column 474   Coefficient 0.60937500
   "01001111", -- Column 475   Coefficient 0.61718750
   "01010000", -- Column 476   Coefficient 0.62500000
   "01010000", -- Column 477   Coefficient 0.62500000
   "01010000", -- Column 478   Coefficient 0.62500000
   "01010000", -- Column 479   Coefficient 0.62500000
   "01010001", -- Column 480   Coefficient 0.63281250
   "01010010", -- Column 481   Coefficient 0.64062500
   "01010011", -- Column 482   Coefficient 0.64843750
   "01010100", -- Column 483   Coefficient 0.65625000
   "01010100", -- Column 484   Coefficient 0.65625000
   "01010100", -- Column 485   Coefficient 0.65625000
   "01010100", -- Column 486   Coefficient 0.65625000
   "01010100", -- Column 487   Coefficient 0.65625000
   "01010110", -- Column 488   Coefficient 0.67187500
   "01010110", -- Column 489   Coefficient 0.67187500
   "01010101", -- Column 490   Coefficient 0.66406250
   "01010101", -- Column 491   Coefficient 0.66406250
   "01010101", -- Column 492   Coefficient 0.66406250
   "01010110", -- Column 493   Coefficient 0.67187500
   "01010110", -- Column 494   Coefficient 0.67187500
   "01010111", -- Column 495   Coefficient 0.67968750
   "01010111", -- Column 496   Coefficient 0.67968750
   "01011000", -- Column 497   Coefficient 0.68750000
   "01011000", -- Column 498   Coefficient 0.68750000
   "01011001", -- Column 499   Coefficient 0.69531250
   "01011001", -- Column 500   Coefficient 0.69531250
   "01011001", -- Column 501   Coefficient 0.69531250
   "01011001", -- Column 502   Coefficient 0.69531250
   "01011010", -- Column 503   Coefficient 0.70312500
   "01011011", -- Column 504   Coefficient 0.71093750
   "01011100", -- Column 505   Coefficient 0.71875000
   "01011100", -- Column 506   Coefficient 0.71875000
   "01011100", -- Column 507   Coefficient 0.71875000
   "01011011", -- Column 508   Coefficient 0.71093750
   "01011100", -- Column 509   Coefficient 0.71875000
   "01011110", -- Column 510   Coefficient 0.73437500
   "01011110", -- Column 511   Coefficient 0.73437500
   "01011110", -- Column 512   Coefficient 0.73437500
   "01011110", -- Column 513   Coefficient 0.73437500
   "01011110", -- Column 514   Coefficient 0.73437500
   "01011111", -- Column 515   Coefficient 0.74218750
   "01100000", -- Column 516   Coefficient 0.75000000
   "01100001", -- Column 517   Coefficient 0.75781250
   "01100001", -- Column 518   Coefficient 0.75781250
   "01100010", -- Column 519   Coefficient 0.76562500
   "01100010", -- Column 520   Coefficient 0.76562500
   "01100010", -- Column 521   Coefficient 0.76562500
   "01100010", -- Column 522   Coefficient 0.76562500
   "01100010", -- Column 523   Coefficient 0.76562500
   "01100011", -- Column 524   Coefficient 0.77343750
   "01100011", -- Column 525   Coefficient 0.77343750
   "01100100", -- Column 526   Coefficient 0.78125000
   "01100100", -- Column 527   Coefficient 0.78125000
   "01100100", -- Column 528   Coefficient 0.78125000
   "01100100", -- Column 529   Coefficient 0.78125000
   "01100100", -- Column 530   Coefficient 0.78125000
   "01100100", -- Column 531   Coefficient 0.78125000
   "01100101", -- Column 532   Coefficient 0.78906250
   "01100101", -- Column 533   Coefficient 0.78906250
   "01100110", -- Column 534   Coefficient 0.79687500
   "01100110", -- Column 535   Coefficient 0.79687500
   "01100110", -- Column 536   Coefficient 0.79687500
   "01100110", -- Column 537   Coefficient 0.79687500
   "01100111", -- Column 538   Coefficient 0.80468750
   "01100111", -- Column 539   Coefficient 0.80468750
   "01100110", -- Column 540   Coefficient 0.79687500
   "01100110", -- Column 541   Coefficient 0.79687500
   "01100110", -- Column 542   Coefficient 0.79687500
   "01100110", -- Column 543   Coefficient 0.79687500
   "01100111", -- Column 544   Coefficient 0.80468750
   "01100111", -- Column 545   Coefficient 0.80468750
   "01100111", -- Column 546   Coefficient 0.80468750
   "01101000", -- Column 547   Coefficient 0.81250000
   "01101000", -- Column 548   Coefficient 0.81250000
   "01101000", -- Column 549   Coefficient 0.81250000
   "01101000", -- Column 550   Coefficient 0.81250000
   "01101000", -- Column 551   Coefficient 0.81250000
   "01101000", -- Column 552   Coefficient 0.81250000
   "01101000", -- Column 553   Coefficient 0.81250000
   "01101000", -- Column 554   Coefficient 0.81250000
   "01101000", -- Column 555   Coefficient 0.81250000
   "01101000", -- Column 556   Coefficient 0.81250000
   "01101000", -- Column 557   Coefficient 0.81250000
   "01100111", -- Column 558   Coefficient 0.80468750
   "01100111", -- Column 559   Coefficient 0.80468750
   "01100111", -- Column 560   Coefficient 0.80468750
   "01100111", -- Column 561   Coefficient 0.80468750
   "01100111", -- Column 562   Coefficient 0.80468750
   "01100110", -- Column 563   Coefficient 0.79687500
   "01100101", -- Column 564   Coefficient 0.78906250
   "01100101", -- Column 565   Coefficient 0.78906250
   "01100110", -- Column 566   Coefficient 0.79687500
   "01100101", -- Column 567   Coefficient 0.78906250
   "01100101", -- Column 568   Coefficient 0.78906250
   "01100101", -- Column 569   Coefficient 0.78906250
   "01100101", -- Column 570   Coefficient 0.78906250
   "01100101", -- Column 571   Coefficient 0.78906250
   "01100100", -- Column 572   Coefficient 0.78125000
   "01100100", -- Column 573   Coefficient 0.78125000
   "01100011", -- Column 574   Coefficient 0.77343750
   "01100011", -- Column 575   Coefficient 0.77343750
   "01100011", -- Column 576   Coefficient 0.77343750
   "01100010", -- Column 577   Coefficient 0.76562500
   "01100001", -- Column 578   Coefficient 0.75781250
   "01100000", -- Column 579   Coefficient 0.75000000
   "01100000", -- Column 580   Coefficient 0.75000000
   "01100000", -- Column 581   Coefficient 0.75000000
   "01011111", -- Column 582   Coefficient 0.74218750
   "01011101", -- Column 583   Coefficient 0.72656250
   "01011101", -- Column 584   Coefficient 0.72656250
   "01011100", -- Column 585   Coefficient 0.71875000
   "01011100", -- Column 586   Coefficient 0.71875000
   "01011010", -- Column 587   Coefficient 0.70312500
   "01011001", -- Column 588   Coefficient 0.69531250
   "01011001", -- Column 589   Coefficient 0.69531250
   "01011001", -- Column 590   Coefficient 0.69531250
   "01010111", -- Column 591   Coefficient 0.67968750
   "01010101", -- Column 592   Coefficient 0.66406250
   "01010100", -- Column 593   Coefficient 0.65625000
   "01010100", -- Column 594   Coefficient 0.65625000
   "01010100", -- Column 595   Coefficient 0.65625000
   "01010010", -- Column 596   Coefficient 0.64062500
   "01010000", -- Column 597   Coefficient 0.62500000
   "01001111", -- Column 598   Coefficient 0.61718750
   "01001111", -- Column 599   Coefficient 0.61718750
   "01001110", -- Column 600   Coefficient 0.60937500
   "01001101", -- Column 601   Coefficient 0.60156250
   "01001100", -- Column 602   Coefficient 0.59375000
   "01001100", -- Column 603   Coefficient 0.59375000
   "01001011", -- Column 604   Coefficient 0.58593750
   "01001010", -- Column 605   Coefficient 0.57812500
   "01001001", -- Column 606   Coefficient 0.57031250
   "01000111", -- Column 607   Coefficient 0.55468750
   "01000101", -- Column 608   Coefficient 0.53906250
   "01000100", -- Column 609   Coefficient 0.53125000
   "01000100", -- Column 610   Coefficient 0.53125000
   "01000100", -- Column 611   Coefficient 0.53125000
   "01000011", -- Column 612   Coefficient 0.52343750
   "01000001", -- Column 613   Coefficient 0.50781250
   "01000000", -- Column 614   Coefficient 0.50000000
   "00111111", -- Column 615   Coefficient 0.49218750
   "00111111", -- Column 616   Coefficient 0.49218750
   "00111110", -- Column 617   Coefficient 0.48437500
   "00111101", -- Column 618   Coefficient 0.47656250
   "00111101", -- Column 619   Coefficient 0.47656250
   "00111101", -- Column 620   Coefficient 0.47656250
   "00111011", -- Column 621   Coefficient 0.46093750
   "00111010", -- Column 622   Coefficient 0.45312500
   "00111001", -- Column 623   Coefficient 0.44531250
   "00111000", -- Column 624   Coefficient 0.43750000
   "00110111", -- Column 625   Coefficient 0.42968750
   "00110111", -- Column 626   Coefficient 0.42968750
   "00110110", -- Column 627   Coefficient 0.42187500
   "00110110", -- Column 628   Coefficient 0.42187500
   "00110110", -- Column 629   Coefficient 0.42187500
   "00110101", -- Column 630   Coefficient 0.41406250
   "00110101", -- Column 631   Coefficient 0.41406250
   "00110100", -- Column 632   Coefficient 0.40625000
   "00110100", -- Column 633   Coefficient 0.40625000
   "00110011", -- Column 634   Coefficient 0.39843750
   "00110011", -- Column 635   Coefficient 0.39843750
   "00110010", -- Column 636   Coefficient 0.39062500
   "00110001", -- Column 637   Coefficient 0.38281250
   "00110000", -- Column 638   Coefficient 0.37500000
   "00110000", -- Column 639   Coefficient 0.37500000
   "00101111", -- Column 640   Coefficient 0.36718750
   "00101110", -- Column 641   Coefficient 0.35937500
   "00101110", -- Column 642   Coefficient 0.35937500
   "00101110", -- Column 643   Coefficient 0.35937500
   "00101110", -- Column 644   Coefficient 0.35937500
   "00101110", -- Column 645   Coefficient 0.35937500
   "00101110", -- Column 646   Coefficient 0.35937500
   "00101101", -- Column 647   Coefficient 0.35156250
   "00101101", -- Column 648   Coefficient 0.35156250
   "00101101", -- Column 649   Coefficient 0.35156250
   "00101101", -- Column 650   Coefficient 0.35156250
   "00101100", -- Column 651   Coefficient 0.34375000
   "00101100", -- Column 652   Coefficient 0.34375000
   "00101011", -- Column 653   Coefficient 0.33593750
   "00101100", -- Column 654   Coefficient 0.34375000
   "00101011", -- Column 655   Coefficient 0.33593750
   "00101011", -- Column 656   Coefficient 0.33593750
   "00101011", -- Column 657   Coefficient 0.33593750
   "00101011", -- Column 658   Coefficient 0.33593750
   "00101010", -- Column 659   Coefficient 0.32812500
   "00101010", -- Column 660   Coefficient 0.32812500
   "00101010", -- Column 661   Coefficient 0.32812500
   "00101010", -- Column 662   Coefficient 0.32812500
   "00101010", -- Column 663   Coefficient 0.32812500
   "00101010", -- Column 664   Coefficient 0.32812500
   "00101001", -- Column 665   Coefficient 0.32031250
   "00101010", -- Column 666   Coefficient 0.32812500
   "00101010", -- Column 667   Coefficient 0.32812500
   "00101010", -- Column 668   Coefficient 0.32812500
   "00101010", -- Column 669   Coefficient 0.32812500
   "00101010", -- Column 670   Coefficient 0.32812500
   "00101010", -- Column 671   Coefficient 0.32812500
   "00101010", -- Column 672   Coefficient 0.32812500
   "00101010", -- Column 673   Coefficient 0.32812500
   "00101010", -- Column 674   Coefficient 0.32812500
   "00101010", -- Column 675   Coefficient 0.32812500
   "00101011", -- Column 676   Coefficient 0.33593750
   "00101010", -- Column 677   Coefficient 0.32812500
   "00101010", -- Column 678   Coefficient 0.32812500
   "00101010", -- Column 679   Coefficient 0.32812500
   "00101011", -- Column 680   Coefficient 0.33593750
   "00101011", -- Column 681   Coefficient 0.33593750
   "00101011", -- Column 682   Coefficient 0.33593750
   "00101010", -- Column 683   Coefficient 0.32812500
   "00101001", -- Column 684   Coefficient 0.32031250
   "00101010", -- Column 685   Coefficient 0.32812500
   "00101011", -- Column 686   Coefficient 0.33593750
   "00101011", -- Column 687   Coefficient 0.33593750
   "00101100", -- Column 688   Coefficient 0.34375000
   "00101011", -- Column 689   Coefficient 0.33593750
   "00101100", -- Column 690   Coefficient 0.34375000
   "00101011", -- Column 691   Coefficient 0.33593750
   "00101011", -- Column 692   Coefficient 0.33593750
   "00101011", -- Column 693   Coefficient 0.33593750
   "00101100", -- Column 694   Coefficient 0.34375000
   "00101100", -- Column 695   Coefficient 0.34375000
   "00101100", -- Column 696   Coefficient 0.34375000
   "00101100", -- Column 697   Coefficient 0.34375000
   "00101100", -- Column 698   Coefficient 0.34375000
   "00101100", -- Column 699   Coefficient 0.34375000
   "00101100", -- Column 700   Coefficient 0.34375000
   "00101100", -- Column 701   Coefficient 0.34375000
   "00101100", -- Column 702   Coefficient 0.34375000
   "00101100", -- Column 703   Coefficient 0.34375000
   "00101101", -- Column 704   Coefficient 0.35156250
   "00101101", -- Column 705   Coefficient 0.35156250
   "00101101", -- Column 706   Coefficient 0.35156250
   "00101100", -- Column 707   Coefficient 0.34375000
   "00101101", -- Column 708   Coefficient 0.35156250
   "00101101", -- Column 709   Coefficient 0.35156250
   "00101101", -- Column 710   Coefficient 0.35156250
   "00101101", -- Column 711   Coefficient 0.35156250
   "00101110", -- Column 712   Coefficient 0.35937500
   "00101110", -- Column 713   Coefficient 0.35937500
   "00101110", -- Column 714   Coefficient 0.35937500
   "00101101", -- Column 715   Coefficient 0.35156250
   "00101101", -- Column 716   Coefficient 0.35156250
   "00101110", -- Column 717   Coefficient 0.35937500
   "00101110", -- Column 718   Coefficient 0.35937500
   "00101101", -- Column 719   Coefficient 0.35156250
   "00101101", -- Column 720   Coefficient 0.35156250
   "00101101", -- Column 721   Coefficient 0.35156250
   "00101110", -- Column 722   Coefficient 0.35937500
   "00101101", -- Column 723   Coefficient 0.35156250
   "00101101", -- Column 724   Coefficient 0.35156250
   "00101100", -- Column 725   Coefficient 0.34375000
   "00101100", -- Column 726   Coefficient 0.34375000
   "00101101", -- Column 727   Coefficient 0.35156250
   "00101110", -- Column 728   Coefficient 0.35937500
   "00101110", -- Column 729   Coefficient 0.35937500
   "00101110", -- Column 730   Coefficient 0.35937500
   "00101110", -- Column 731   Coefficient 0.35937500
   "00101101", -- Column 732   Coefficient 0.35156250
   "00101101", -- Column 733   Coefficient 0.35156250
   "00101101", -- Column 734   Coefficient 0.35156250
   "00101110", -- Column 735   Coefficient 0.35937500
   "00101111", -- Column 736   Coefficient 0.36718750
   "00101110", -- Column 737   Coefficient 0.35937500
   "00101110", -- Column 738   Coefficient 0.35937500
   "00101110", -- Column 739   Coefficient 0.35937500
   "00101110", -- Column 740   Coefficient 0.35937500
   "00101110", -- Column 741   Coefficient 0.35937500
   "00101110", -- Column 742   Coefficient 0.35937500
   "00101101", -- Column 743   Coefficient 0.35156250
   "00101101", -- Column 744   Coefficient 0.35156250
   "00101101", -- Column 745   Coefficient 0.35156250
   "00101101", -- Column 746   Coefficient 0.35156250
   "00101101", -- Column 747   Coefficient 0.35156250
   "00101110", -- Column 748   Coefficient 0.35937500
   "00101110", -- Column 749   Coefficient 0.35937500
   "00101110", -- Column 750   Coefficient 0.35937500
   "00101110", -- Column 751   Coefficient 0.35937500
   "00101110", -- Column 752   Coefficient 0.35937500
   "00101110", -- Column 753   Coefficient 0.35937500
   "00101101", -- Column 754   Coefficient 0.35156250
   "00101101", -- Column 755   Coefficient 0.35156250
   "00101110", -- Column 756   Coefficient 0.35937500
   "00101110", -- Column 757   Coefficient 0.35937500
   "00101110", -- Column 758   Coefficient 0.35937500
   "00101101", -- Column 759   Coefficient 0.35156250
   "00101101", -- Column 760   Coefficient 0.35156250
   "00101110", -- Column 761   Coefficient 0.35937500
   "00101110", -- Column 762   Coefficient 0.35937500
   "00101110", -- Column 763   Coefficient 0.35937500
   "00101110", -- Column 764   Coefficient 0.35937500
   "00101101", -- Column 765   Coefficient 0.35156250
   "00101100", -- Column 766   Coefficient 0.34375000
   "00101100", -- Column 767   Coefficient 0.34375000
   "00101101", -- Column 768   Coefficient 0.35156250
   "00101110", -- Column 769   Coefficient 0.35937500
   "00101110", -- Column 770   Coefficient 0.35937500
   "00101101", -- Column 771   Coefficient 0.35156250
   "00101101", -- Column 772   Coefficient 0.35156250
   "00101101", -- Column 773   Coefficient 0.35156250
   "00101101", -- Column 774   Coefficient 0.35156250
   "00101100", -- Column 775   Coefficient 0.34375000
   "00101100", -- Column 776   Coefficient 0.34375000
   "00101100", -- Column 777   Coefficient 0.34375000
   "00101101", -- Column 778   Coefficient 0.35156250
   "00101100", -- Column 779   Coefficient 0.34375000
   "00101100", -- Column 780   Coefficient 0.34375000
   "00101100", -- Column 781   Coefficient 0.34375000
   "00101100", -- Column 782   Coefficient 0.34375000
   "00101100", -- Column 783   Coefficient 0.34375000
   "00101011", -- Column 784   Coefficient 0.33593750
   "00101011", -- Column 785   Coefficient 0.33593750
   "00101011", -- Column 786   Coefficient 0.33593750
   "00101011", -- Column 787   Coefficient 0.33593750
   "00101011", -- Column 788   Coefficient 0.33593750
   "00101011", -- Column 789   Coefficient 0.33593750
   "00101011", -- Column 790   Coefficient 0.33593750
   "00101011", -- Column 791   Coefficient 0.33593750
   "00101011", -- Column 792   Coefficient 0.33593750
   "00101011", -- Column 793   Coefficient 0.33593750
   "00101010", -- Column 794   Coefficient 0.32812500
   "00101010", -- Column 795   Coefficient 0.32812500
   "00101010", -- Column 796   Coefficient 0.32812500
   "00101010", -- Column 797   Coefficient 0.32812500
   "00101010", -- Column 798   Coefficient 0.32812500
   "00101001", -- Column 799   Coefficient 0.32031250
   "00101001", -- Column 800   Coefficient 0.32031250
   "00101010", -- Column 801   Coefficient 0.32812500
   "00101001", -- Column 802   Coefficient 0.32031250
   "00101001", -- Column 803   Coefficient 0.32031250
   "00101001", -- Column 804   Coefficient 0.32031250
   "00101001", -- Column 805   Coefficient 0.32031250
   "00101001", -- Column 806   Coefficient 0.32031250
   "00101000", -- Column 807   Coefficient 0.31250000
   "00101000", -- Column 808   Coefficient 0.31250000
   "00101000", -- Column 809   Coefficient 0.31250000
   "00101000", -- Column 810   Coefficient 0.31250000
   "00101000", -- Column 811   Coefficient 0.31250000
   "00101000", -- Column 812   Coefficient 0.31250000
   "00101001", -- Column 813   Coefficient 0.32031250
   "00101001", -- Column 814   Coefficient 0.32031250
   "00101001", -- Column 815   Coefficient 0.32031250
   "00101001", -- Column 816   Coefficient 0.32031250
   "00101001", -- Column 817   Coefficient 0.32031250
   "00101000", -- Column 818   Coefficient 0.31250000
   "00101000", -- Column 819   Coefficient 0.31250000
   "00100111", -- Column 820   Coefficient 0.30468750
   "00100111", -- Column 821   Coefficient 0.30468750
   "00101000", -- Column 822   Coefficient 0.31250000
   "00101000", -- Column 823   Coefficient 0.31250000
   "00101000", -- Column 824   Coefficient 0.31250000
   "00100111", -- Column 825   Coefficient 0.30468750
   "00100110", -- Column 826   Coefficient 0.29687500
   "00100110", -- Column 827   Coefficient 0.29687500
   "00100110", -- Column 828   Coefficient 0.29687500
   "00100111", -- Column 829   Coefficient 0.30468750
   "00100111", -- Column 830   Coefficient 0.30468750
   "00100111", -- Column 831   Coefficient 0.30468750
   "00100111", -- Column 832   Coefficient 0.30468750
   "00100111", -- Column 833   Coefficient 0.30468750
   "00100110", -- Column 834   Coefficient 0.29687500
   "00100110", -- Column 835   Coefficient 0.29687500
   "00100111", -- Column 836   Coefficient 0.30468750
   "00100111", -- Column 837   Coefficient 0.30468750
   "00100111", -- Column 838   Coefficient 0.30468750
   "00100110", -- Column 839   Coefficient 0.29687500
   "00100110", -- Column 840   Coefficient 0.29687500
   "00100110", -- Column 841   Coefficient 0.29687500
   "00100110", -- Column 842   Coefficient 0.29687500
   "00100101", -- Column 843   Coefficient 0.28906250
   "00100101", -- Column 844   Coefficient 0.28906250
   "00100110", -- Column 845   Coefficient 0.29687500
   "00100110", -- Column 846   Coefficient 0.29687500
   "00100110", -- Column 847   Coefficient 0.29687500
   "00100110", -- Column 848   Coefficient 0.29687500
   "00100110", -- Column 849   Coefficient 0.29687500
   "00100110", -- Column 850   Coefficient 0.29687500
   "00100110", -- Column 851   Coefficient 0.29687500
   "00100101", -- Column 852   Coefficient 0.28906250
   "00100101", -- Column 853   Coefficient 0.28906250
   "00100101", -- Column 854   Coefficient 0.28906250
   "00100101", -- Column 855   Coefficient 0.28906250
   "00100101", -- Column 856   Coefficient 0.28906250
   "00100100", -- Column 857   Coefficient 0.28125000
   "00100100", -- Column 858   Coefficient 0.28125000
   "00100100", -- Column 859   Coefficient 0.28125000
   "00100101", -- Column 860   Coefficient 0.28906250
   "00100101", -- Column 861   Coefficient 0.28906250
   "00100101", -- Column 862   Coefficient 0.28906250
   "00100101", -- Column 863   Coefficient 0.28906250
   "00100100", -- Column 864   Coefficient 0.28125000
   "00100101", -- Column 865   Coefficient 0.28906250
   "00100101", -- Column 866   Coefficient 0.28906250
   "00100101", -- Column 867   Coefficient 0.28906250
   "00100101", -- Column 868   Coefficient 0.28906250
   "00100110", -- Column 869   Coefficient 0.29687500
   "00100110", -- Column 870   Coefficient 0.29687500
   "00100101", -- Column 871   Coefficient 0.28906250
   "00100100", -- Column 872   Coefficient 0.28125000
   "00100100", -- Column 873   Coefficient 0.28125000
   "00100100", -- Column 874   Coefficient 0.28125000
   "00100100", -- Column 875   Coefficient 0.28125000
   "00100100", -- Column 876   Coefficient 0.28125000
   "00100100", -- Column 877   Coefficient 0.28125000
   "00100100", -- Column 878   Coefficient 0.28125000
   "00100100", -- Column 879   Coefficient 0.28125000
   "00100011", -- Column 880   Coefficient 0.27343750
   "00100011", -- Column 881   Coefficient 0.27343750
   "00100100", -- Column 882   Coefficient 0.28125000
   "00100011", -- Column 883   Coefficient 0.27343750
   "00100011", -- Column 884   Coefficient 0.27343750
   "00100011", -- Column 885   Coefficient 0.27343750
   "00100100", -- Column 886   Coefficient 0.28125000
   "00100100", -- Column 887   Coefficient 0.28125000
   "00100100", -- Column 888   Coefficient 0.28125000
   "00100100", -- Column 889   Coefficient 0.28125000
   "00100100", -- Column 890   Coefficient 0.28125000
   "00100101", -- Column 891   Coefficient 0.28906250
   "00100101", -- Column 892   Coefficient 0.28906250
   "00100011", -- Column 893   Coefficient 0.27343750
   "00100011", -- Column 894   Coefficient 0.27343750
   "00100011", -- Column 895   Coefficient 0.27343750
   "00100011", -- Column 896   Coefficient 0.27343750
   "00100011", -- Column 897   Coefficient 0.27343750
   "00100011", -- Column 898   Coefficient 0.27343750
   "00100011", -- Column 899   Coefficient 0.27343750
   "00100100", -- Column 900   Coefficient 0.28125000
   "00100100", -- Column 901   Coefficient 0.28125000
   "00100100", -- Column 902   Coefficient 0.28125000
   "00100011", -- Column 903   Coefficient 0.27343750
   "00100011", -- Column 904   Coefficient 0.27343750
   "00100011", -- Column 905   Coefficient 0.27343750
   "00100010", -- Column 906   Coefficient 0.26562500
   "00100010", -- Column 907   Coefficient 0.26562500
   "00100011", -- Column 908   Coefficient 0.27343750
   "00100011", -- Column 909   Coefficient 0.27343750
   "00100100", -- Column 910   Coefficient 0.28125000
   "00100011", -- Column 911   Coefficient 0.27343750
   "00100100", -- Column 912   Coefficient 0.28125000
   "00100100", -- Column 913   Coefficient 0.28125000
   "00100100", -- Column 914   Coefficient 0.28125000
   "00100011", -- Column 915   Coefficient 0.27343750
   "00100100", -- Column 916   Coefficient 0.28125000
   "00100100", -- Column 917   Coefficient 0.28125000
   "00100100", -- Column 918   Coefficient 0.28125000
   "00100011", -- Column 919   Coefficient 0.27343750
   "00100010", -- Column 920   Coefficient 0.26562500
   "00100010", -- Column 921   Coefficient 0.26562500
   "00100010", -- Column 922   Coefficient 0.26562500
   "00100011", -- Column 923   Coefficient 0.27343750
   "00100011", -- Column 924   Coefficient 0.27343750
   "00100010", -- Column 925   Coefficient 0.26562500
   "00100010", -- Column 926   Coefficient 0.26562500
   "00100011", -- Column 927   Coefficient 0.27343750
   "00100011", -- Column 928   Coefficient 0.27343750
   "00100011", -- Column 929   Coefficient 0.27343750
   "00100011", -- Column 930   Coefficient 0.27343750
   "00100010", -- Column 931   Coefficient 0.26562500
   "00100010", -- Column 932   Coefficient 0.26562500
   "00100011", -- Column 933   Coefficient 0.27343750
   "00100011", -- Column 934   Coefficient 0.27343750
   "00100011", -- Column 935   Coefficient 0.27343750
   "00100011", -- Column 936   Coefficient 0.27343750
   "00100011", -- Column 937   Coefficient 0.27343750
   "00100010", -- Column 938   Coefficient 0.26562500
   "00100010", -- Column 939   Coefficient 0.26562500
   "00100010", -- Column 940   Coefficient 0.26562500
   "00100010", -- Column 941   Coefficient 0.26562500
   "00100010", -- Column 942   Coefficient 0.26562500
   "00100010", -- Column 943   Coefficient 0.26562500
   "00100010", -- Column 944   Coefficient 0.26562500
   "00100011", -- Column 945   Coefficient 0.27343750
   "00100011", -- Column 946   Coefficient 0.27343750
   "00100011", -- Column 947   Coefficient 0.27343750
   "00100011", -- Column 948   Coefficient 0.27343750
   "00100011", -- Column 949   Coefficient 0.27343750
   "00100011", -- Column 950   Coefficient 0.27343750
   "00100100", -- Column 951   Coefficient 0.28125000
   "00100100", -- Column 952   Coefficient 0.28125000
   "00100100", -- Column 953   Coefficient 0.28125000
   "00100100", -- Column 954   Coefficient 0.28125000
   "00100100", -- Column 955   Coefficient 0.28125000
   "00100100", -- Column 956   Coefficient 0.28125000
   "00100011", -- Column 957   Coefficient 0.27343750
   "00100011", -- Column 958   Coefficient 0.27343750
   "00100100", -- Column 959   Coefficient 0.28125000
   "00100100", -- Column 960   Coefficient 0.28125000
   "00100101", -- Column 961   Coefficient 0.28906250
   "00100101", -- Column 962   Coefficient 0.28906250
   "00100110", -- Column 963   Coefficient 0.29687500
   "00100110", -- Column 964   Coefficient 0.29687500
   "00100110", -- Column 965   Coefficient 0.29687500
   "00100101", -- Column 966   Coefficient 0.28906250
   "00100110", -- Column 967   Coefficient 0.29687500
   "00100110", -- Column 968   Coefficient 0.29687500
   "00100111", -- Column 969   Coefficient 0.30468750
   "00100111", -- Column 970   Coefficient 0.30468750
   "00100111", -- Column 971   Coefficient 0.30468750
   "00101000", -- Column 972   Coefficient 0.31250000
   "00101001", -- Column 973   Coefficient 0.32031250
   "00101001", -- Column 974   Coefficient 0.32031250
   "00101000", -- Column 975   Coefficient 0.31250000
   "00101000", -- Column 976   Coefficient 0.31250000
   "00101001", -- Column 977   Coefficient 0.32031250
   "00101010", -- Column 978   Coefficient 0.32812500
   "00101010", -- Column 979   Coefficient 0.32812500
   "00101011", -- Column 980   Coefficient 0.33593750
   "00101011", -- Column 981   Coefficient 0.33593750
   "00101100", -- Column 982   Coefficient 0.34375000
   "00101100", -- Column 983   Coefficient 0.34375000
   "00101100", -- Column 984   Coefficient 0.34375000
   "00101100", -- Column 985   Coefficient 0.34375000
   "00101100", -- Column 986   Coefficient 0.34375000
   "00101100", -- Column 987   Coefficient 0.34375000
   "00101101", -- Column 988   Coefficient 0.35156250
   "00101101", -- Column 989   Coefficient 0.35156250
   "00101101", -- Column 990   Coefficient 0.35156250
   "00101101", -- Column 991   Coefficient 0.35156250
   "00101101", -- Column 992   Coefficient 0.35156250
   "00101101", -- Column 993   Coefficient 0.35156250
   "00101101", -- Column 994   Coefficient 0.35156250
   "00101100", -- Column 995   Coefficient 0.34375000
   "00101011", -- Column 996   Coefficient 0.33593750
   "00101011", -- Column 997   Coefficient 0.33593750
   "00101011", -- Column 998   Coefficient 0.33593750
   "00101011", -- Column 999   Coefficient 0.33593750
   "00101100", -- Column 1000   Coefficient 0.34375000
   "00101101", -- Column 1001   Coefficient 0.35156250
   "00101110", -- Column 1002   Coefficient 0.35937500
   "00101101", -- Column 1003   Coefficient 0.35156250
   "00101101", -- Column 1004   Coefficient 0.35156250
   "00101100", -- Column 1005   Coefficient 0.34375000
   "00101101", -- Column 1006   Coefficient 0.35156250
   "00101101", -- Column 1007   Coefficient 0.35156250
   "00101101", -- Column 1008   Coefficient 0.35156250
   "00101101", -- Column 1009   Coefficient 0.35156250
   "00101101", -- Column 1010   Coefficient 0.35156250
   "00101101", -- Column 1011   Coefficient 0.35156250
   "00101110", -- Column 1012   Coefficient 0.35937500
   "00101101", -- Column 1013   Coefficient 0.35156250
   "00101100", -- Column 1014   Coefficient 0.34375000
   "00101100", -- Column 1015   Coefficient 0.34375000
   "00101101", -- Column 1016   Coefficient 0.35156250
   "00101110", -- Column 1017   Coefficient 0.35937500
   "00101110", -- Column 1018   Coefficient 0.35937500
   "00101101", -- Column 1019   Coefficient 0.35156250
   "00101101", -- Column 1020   Coefficient 0.35156250
   "00101100", -- Column 1021   Coefficient 0.34375000
   "00101100", -- Column 1022   Coefficient 0.34375000
   "00101011", -- Column 1023   Coefficient 0.33593750
   "00101011" -- Column 1024   Coefficient 0.33593750
);
begin
	process(clk)
	begin
	if(rising_edge(CLK)) then
		A <= rom(to_integer(unsigned(I)));
	end if;
	end process;
end ROM;
