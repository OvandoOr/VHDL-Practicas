library ieee; 
use ieee.std_logic_1164.all;	
use ieee.numeric_std.all;
entity Rom_Histograma_sine is
	generic(
	n: 	integer:= 12;		-- No. de bits informacion
	m:	integer:= 9 		-- No. de bits para datos
	); 
	port 
	(
		CLK		: in std_logic;
		addr	: in std_logic_vector (m-1 downto 0);
		q		: out std_logic_vector((n -1) downto 0)
	);
end Rom_Histograma_sine;
architecture rtl of Rom_Histograma_sine is
	subtype word_t is std_logic_vector((n-1) downto 0);
	type memory_t is array(0 to (2**m)-1 ) of word_t;
	function init_rom
		return memory_t is 
		variable tmp : memory_t :=(
	 "110001110001",  	 --  3185 	 0 
	 "110011001100",  	 --  3276 	 1 
	 "110100100110",  	 --  3366 	 2 
	 "110101111110",  	 --  3454 	 3 
	 "110111010011",  	 --  3539 	 4 
	 "111000100101",  	 --  3621 	 5 
	 "111001110011",  	 --  3699 	 6 
	 "111010111011",  	 --  3771 	 7 
	 "111011111110",  	 --  3838 	 8 
	 "111100111010",  	 --  3898 	 9 
	 "111101101111",  	 --  3951 	 10 
	 "111110011100",  	 --  3996 	 11 
	 "111111000001",  	 --  4033 	 12 
	 "111111011110",  	 --  4062 	 13 
	 "111111110010",  	 --  4082 	 14 
	 "111111111101",  	 --  4093 	 15 
	 "111111111111",  	 --  4095 	 16 
	 "111111110111",  	 --  4087 	 17 
	 "111111100111",  	 --  4071 	 18 
	 "111111001110",  	 --  4046 	 19 
	 "111110101100",  	 --  4012 	 20 
	 "111110000011",  	 --  3971 	 21 
	 "111101010001",  	 --  3921 	 22 
	 "111100011000",  	 --  3864 	 23 
	 "111011011000",  	 --  3800 	 24 
	 "111010010010",  	 --  3730 	 25 
	 "111001000110",  	 --  3654 	 26 
	 "110111110110",  	 --  3574 	 27 
	 "110110100010",  	 --  3490 	 28 
	 "110101001011",  	 --  3403 	 29 
	 "110011110001",  	 --  3313 	 30 
	 "110010010111",  	 --  3223 	 31 
	 "110000111100",  	 --  3132 	 32 
	 "101111100001",  	 --  3041 	 33 
	 "101110001000",  	 --  2952 	 34 
	 "101100110010",  	 --  2866 	 35 
	 "101011011110",  	 --  2782 	 36 
	 "101010001111",  	 --  2703 	 37 
	 "101001000100",  	 --  2628 	 38 
	 "100111111111",  	 --  2559 	 39 
	 "100111000000",  	 --  2496 	 40 
	 "100110001000",  	 --  2440 	 41 
	 "100101011000",  	 --  2392 	 42 
	 "100100101111",  	 --  2351 	 43 
	 "100100001111",  	 --  2319 	 44 
	 "100011110111",  	 --  2295 	 45 
	 "100011101001",  	 --  2281 	 46 
	 "100011100011",  	 --  2275 	 47 
	 "100011100110",  	 --  2278 	 48 
	 "100011110011",  	 --  2291 	 49 
	 "100100001000",  	 --  2312 	 50 
	 "100100100111",  	 --  2343 	 51 
	 "100101001101",  	 --  2381 	 52 
	 "100101111100",  	 --  2428 	 53 
	 "100110110010",  	 --  2482 	 54 
	 "100111101111",  	 --  2543 	 55 
	 "101000110011",  	 --  2611 	 56 
	 "101001111100",  	 --  2684 	 57 
	 "101011001010",  	 --  2762 	 58 
	 "101100011101",  	 --  2845 	 59 
	 "101101110011",  	 --  2931 	 60 
	 "101111001011",  	 --  3019 	 61 
	 "110000100101",  	 --  3109 	 62 
	 "110010000000",  	 --  3200 	 63 
	 "110011011011",  	 --  3291 	 64 
	 "110100110101",  	 --  3381 	 65 
	 "110110001101",  	 --  3469 	 66 
	 "110111100001",  	 --  3553 	 67 
	 "111000110011",  	 --  3635 	 68 
	 "111001111111",  	 --  3711 	 69 
	 "111011000111",  	 --  3783 	 70 
	 "111100001000",  	 --  3848 	 71 
	 "111101000011",  	 --  3907 	 72 
	 "111101110111",  	 --  3959 	 73 
	 "111110100011",  	 --  4003 	 74 
	 "111111000111",  	 --  4039 	 75 
	 "111111100010",  	 --  4066 	 76 
	 "111111110100",  	 --  4084 	 77 
	 "111111111110",  	 --  4094 	 78 
	 "111111111110",  	 --  4094 	 79 
	 "111111110101",  	 --  4085 	 80 
	 "111111100100",  	 --  4068 	 81 
	 "111111001001",  	 --  4041 	 82 
	 "111110100110",  	 --  4006 	 83 
	 "111101111011",  	 --  3963 	 84 
	 "111101001000",  	 --  3912 	 85 
	 "111100001101",  	 --  3853 	 86 
	 "111011001100",  	 --  3788 	 87 
	 "111010000101",  	 --  3717 	 88 
	 "111000111001",  	 --  3641 	 89 
	 "110111101000",  	 --  3560 	 90 
	 "110110010011",  	 --  3475 	 91 
	 "110100111100",  	 --  3388 	 92 
	 "110011100010",  	 --  3298 	 93 
	 "110010001000",  	 --  3208 	 94 
	 "110000101101",  	 --  3117 	 95 
	 "101111010010",  	 --  3026 	 96 
	 "101101111010",  	 --  2938 	 97 
	 "101100100100",  	 --  2852 	 98 
	 "101011010001",  	 --  2769 	 99 
	 "101010000010",  	 --  2690 	 100 
	 "101000111000",  	 --  2616 	 101 
	 "100111110100",  	 --  2548 	 102 
	 "100110110110",  	 --  2486 	 103 
	 "100110000000",  	 --  2432 	 104 
	 "100101010000",  	 --  2384 	 105 
	 "100100101001",  	 --  2345 	 106 
	 "100100001010",  	 --  2314 	 107 
	 "100011110100",  	 --  2292 	 108 
	 "100011100111",  	 --  2279 	 109 
	 "100011100011",  	 --  2275 	 110 
	 "100011101000",  	 --  2280 	 111 
	 "100011110110",  	 --  2294 	 112 
	 "100100001101",  	 --  2317 	 113 
	 "100100101100",  	 --  2348 	 114 
	 "100101010100",  	 --  2388 	 115 
	 "100110000100",  	 --  2436 	 116 
	 "100110111100",  	 --  2492 	 117 
	 "100111111010",  	 --  2554 	 118 
	 "101000111110",  	 --  2622 	 119 
	 "101010001001",  	 --  2697 	 120 
	 "101011011000",  	 --  2776 	 121 
	 "101100101011",  	 --  2859 	 122 
	 "101110000001",  	 --  2945 	 123 
	 "101111011010",  	 --  3034 	 124 
	 "110000110101",  	 --  3125 	 125 
	 "110010010000",  	 --  3216 	 126 
	 "110011101010",  	 --  3306 	 127 
	 "110101000100",  	 --  3396 	 128 
	 "110110011011",  	 --  3483 	 129 
	 "110111101111",  	 --  3567 	 130 
	 "111001000000",  	 --  3648 	 131 
	 "111010001100",  	 --  3724 	 132 
	 "111011010010",  	 --  3794 	 133 
	 "111100010011",  	 --  3859 	 134 
	 "111101001100",  	 --  3916 	 135 
	 "111101111111",  	 --  3967 	 136 
	 "111110101001",  	 --  4009 	 137 
	 "111111001100",  	 --  4044 	 138 
	 "111111100110",  	 --  4070 	 139 
	 "111111110110",  	 --  4086 	 140 
	 "111111111110",  	 --  4094 	 141 
	 "111111111101",  	 --  4093 	 142 
	 "111111110011",  	 --  4083 	 143 
	 "111111100000",  	 --  4064 	 144 
	 "111111000100",  	 --  4036 	 145 
	 "111110011111",  	 --  3999 	 146 
	 "111101110011",  	 --  3955 	 147 
	 "111100111110",  	 --  3902 	 148 
	 "111100000011",  	 --  3843 	 149 
	 "111011000001",  	 --  3777 	 150 
	 "111001111001",  	 --  3705 	 151 
	 "111000101100",  	 --  3628 	 152 
	 "110111011010",  	 --  3546 	 153 
	 "110110000101",  	 --  3461 	 154 
	 "110100101101",  	 --  3373 	 155 
	 "110011010011",  	 --  3283 	 156 
	 "110001111000",  	 --  3192 	 157 
	 "110000011101",  	 --  3101 	 158 
	 "101111000011",  	 --  3011 	 159 
	 "101101101011",  	 --  2923 	 160 
	 "101100010101",  	 --  2837 	 161 
	 "101011000011",  	 --  2755 	 162 
	 "101001110101",  	 --  2677 	 163 
	 "101000101100",  	 --  2604 	 164 
	 "100111101001",  	 --  2537 	 165 
	 "100110101101",  	 --  2477 	 166 
	 "100101110111",  	 --  2423 	 167 
	 "100101001001",  	 --  2377 	 168 
	 "100100100011",  	 --  2339 	 169 
	 "100100000110",  	 --  2310 	 170 
	 "100011110010",  	 --  2290 	 171 
	 "100011100110",  	 --  2278 	 172 
	 "100011100011",  	 --  2275 	 173 
	 "100011101010",  	 --  2282 	 174 
	 "100011111001",  	 --  2297 	 175 
	 "100100010010",  	 --  2322 	 176 
	 "100100110011",  	 --  2355 	 177 
	 "100101011100",  	 --  2396 	 178 
	 "100110001101",  	 --  2445 	 179 
	 "100111000110",  	 --  2502 	 180 
	 "101000000101",  	 --  2565 	 181 
	 "101001001011",  	 --  2635 	 182 
	 "101010010110",  	 --  2710 	 183 
	 "101011100110",  	 --  2790 	 184 
	 "101100111001",  	 --  2873 	 185 
	 "101110010000",  	 --  2960 	 186 
	 "101111101001",  	 --  3049 	 187 
	 "110001000100",  	 --  3140 	 188 
	 "110010011111",  	 --  3231 	 189 
	 "110011111001",  	 --  3321 	 190 
	 "110101010011",  	 --  3411 	 191 
	 "110110101001",  	 --  3497 	 192 
	 "110111111101",  	 --  3581 	 193 
	 "111001001101",  	 --  3661 	 194 
	 "111010011000",  	 --  3736 	 195 
	 "111011011110",  	 --  3806 	 196 
	 "111100011101",  	 --  3869 	 197 
	 "111101010101",  	 --  3925 	 198 
	 "111110000111",  	 --  3975 	 199 
	 "111110110000",  	 --  4016 	 200 
	 "111111010001",  	 --  4049 	 201 
	 "111111101001",  	 --  4073 	 202 
	 "111111111000",  	 --  4088 	 203 
	 "111111111111",  	 --  4095 	 204 
	 "111111111100",  	 --  4092 	 205 
	 "111111110000",  	 --  4080 	 206 
	 "111111011100",  	 --  4060 	 207 
	 "111110111110",  	 --  4030 	 208 
	 "111110011000",  	 --  3992 	 209 
	 "111101101010",  	 --  3946 	 210 
	 "111100110101",  	 --  3893 	 211 
	 "111011111000",  	 --  3832 	 212 
	 "111010110101",  	 --  3765 	 213 
	 "111001101100",  	 --  3692 	 214 
	 "111000011110",  	 --  3614 	 215 
	 "110111001100",  	 --  3532 	 216 
	 "110101110110",  	 --  3446 	 217 
	 "110100011110",  	 --  3358 	 218 
	 "110011000100",  	 --  3268 	 219 
	 "110001101001",  	 --  3177 	 220 
	 "110000001110",  	 --  3086 	 221 
	 "101110110100",  	 --  2996 	 222 
	 "101101011100",  	 --  2908 	 223 
	 "101100000111",  	 --  2823 	 224 
	 "101010110110",  	 --  2742 	 225 
	 "101001101001",  	 --  2665 	 226 
	 "101000100001",  	 --  2593 	 227 
	 "100111011111",  	 --  2527 	 228 
	 "100110100011",  	 --  2467 	 229 
	 "100101101111",  	 --  2415 	 230 
	 "100101000010",  	 --  2370 	 231 
	 "100100011110",  	 --  2334 	 232 
	 "100100000010",  	 --  2306 	 233 
	 "100011101111",  	 --  2287 	 234 
	 "100011100101",  	 --  2277 	 235 
	 "100011100100",  	 --  2276 	 236 
	 "100011101100",  	 --  2284 	 237 
	 "100011111101",  	 --  2301 	 238 
	 "100100010111",  	 --  2327 	 239 
	 "100100111001",  	 --  2361 	 240 
	 "100101100100",  	 --  2404 	 241 
	 "100110010110",  	 --  2454 	 242 
	 "100111010000",  	 --  2512 	 243 
	 "101000010000",  	 --  2576 	 244 
	 "101001010111",  	 --  2647 	 245 
	 "101010100011",  	 --  2723 	 246 
	 "101011110011",  	 --  2803 	 247 
	 "101101001000",  	 --  2888 	 248 
	 "101110011111",  	 --  2975 	 249 
	 "101111111001",  	 --  3065 	 250 
	 "110001010011",  	 --  3155 	 251 
	 "110010101110",  	 --  3246 	 252 
	 "110100001000",  	 --  3336 	 253 
	 "110101100001",  	 --  3425 	 254 
	 "110110111000",  	 --  3512 	 255 
	 "111000001011",  	 --  3595 	 256 
	 "111001011010",  	 --  3674 	 257 
	 "111010100100",  	 --  3748 	 258 
	 "111011101001",  	 --  3817 	 259 
	 "111100100111",  	 --  3879 	 260 
	 "111101011110",  	 --  3934 	 261 
	 "111110001110",  	 --  3982 	 262 
	 "111110110110",  	 --  4022 	 263 
	 "111111010101",  	 --  4053 	 264 
	 "111111101100",  	 --  4076 	 265 
	 "111111111010",  	 --  4090 	 266 
	 "111111111111",  	 --  4095 	 267 
	 "111111111011",  	 --  4091 	 268 
	 "111111101101",  	 --  4077 	 269 
	 "111111010111",  	 --  4055 	 270 
	 "111110111000",  	 --  4024 	 271 
	 "111110010001",  	 --  3985 	 272 
	 "111101100010",  	 --  3938 	 273 
	 "111100101011",  	 --  3883 	 274 
	 "111011101101",  	 --  3821 	 275 
	 "111010101001",  	 --  3753 	 276 
	 "111001011111",  	 --  3679 	 277 
	 "111000010001",  	 --  3601 	 278 
	 "110110111110",  	 --  3518 	 279 
	 "110101101000",  	 --  3432 	 280 
	 "110100001111",  	 --  3343 	 281 
	 "110010110101",  	 --  3253 	 282 
	 "110001011010",  	 --  3162 	 283 
	 "101111111111",  	 --  3071 	 284 
	 "101110100101",  	 --  2981 	 285 
	 "101101001110",  	 --  2894 	 286 
	 "101011111001",  	 --  2809 	 287 
	 "101010101000",  	 --  2728 	 288 
	 "101001011100",  	 --  2652 	 289 
	 "101000010101",  	 --  2581 	 290 
	 "100111010100",  	 --  2516 	 291 
	 "100110011010",  	 --  2458 	 292 
	 "100101100111",  	 --  2407 	 293 
	 "100100111100",  	 --  2364 	 294 
	 "100100011001",  	 --  2329 	 295 
	 "100011111110",  	 --  2302 	 296 
	 "100011101101",  	 --  2285 	 297 
	 "100011100100",  	 --  2276 	 298 
	 "100011100100",  	 --  2276 	 299 
	 "100011101110",  	 --  2286 	 300 
	 "100100000000",  	 --  2304 	 301 
	 "100100011100",  	 --  2332 	 302 
	 "100101000000",  	 --  2368 	 303 
	 "100101101100",  	 --  2412 	 304 
	 "100110011111",  	 --  2463 	 305 
	 "100111011010",  	 --  2522 	 306 
	 "101000011100",  	 --  2588 	 307 
	 "101001100011",  	 --  2659 	 308 
	 "101010110000",  	 --  2736 	 309 
	 "101100000001",  	 --  2817 	 310 
	 "101101010110",  	 --  2902 	 311 
	 "101110101110",  	 --  2990 	 312 
	 "110000001000",  	 --  3080 	 313 
	 "110001100011",  	 --  3171 	 314 
	 "110010111101",  	 --  3261 	 315 
	 "110100011000",  	 --  3352 	 316 
	 "110101110000",  	 --  3440 	 317 
	 "110111000110",  	 --  3526 	 318 
	 "111000011001",  	 --  3609 	 319 
	 "111001100111",  	 --  3687 	 320 
	 "111010110000",  	 --  3760 	 321 
	 "111011110100",  	 --  3828 	 322 
	 "111100110001",  	 --  3889 	 323 
	 "111101100111",  	 --  3943 	 324 
	 "111110010101",  	 --  3989 	 325 
	 "111110111100",  	 --  4028 	 326 
	 "111111011010",  	 --  4058 	 327 
	 "111111101111",  	 --  4079 	 328 
	 "111111111100",  	 --  4092 	 329 
	 "111111111111",  	 --  4095 	 330 
	 "111111111001",  	 --  4089 	 331 
	 "111111101010",  	 --  4074 	 332 
	 "111111010011",  	 --  4051 	 333 
	 "111110110010",  	 --  4018 	 334 
	 "111110001010",  	 --  3978 	 335 
	 "111101011001",  	 --  3929 	 336 
	 "111100100001",  	 --  3873 	 337 
	 "111011100010",  	 --  3810 	 338 
	 "111010011101",  	 --  3741 	 339 
	 "111001010010",  	 --  3666 	 340 
	 "111000000011",  	 --  3587 	 341 
	 "110110101111",  	 --  3503 	 342 
	 "110101011001",  	 --  3417 	 343 
	 "110100000000",  	 --  3328 	 344 
	 "110010100101",  	 --  3237 	 345 
	 "110001001010",  	 --  3146 	 346 
	 "101111110000",  	 --  3056 	 347 
	 "101110010110",  	 --  2966 	 348 
	 "101100111111",  	 --  2879 	 349 
	 "101011101011",  	 --  2795 	 350 
	 "101010011011",  	 --  2715 	 351 
	 "101001010000",  	 --  2640 	 352 
	 "101000001010",  	 --  2570 	 353 
	 "100111001010",  	 --  2506 	 354 
	 "100110010001",  	 --  2449 	 355 
	 "100101011111",  	 --  2399 	 356 
	 "100100110101",  	 --  2357 	 357 
	 "100100010100",  	 --  2324 	 358 
	 "100011111011",  	 --  2299 	 359 
	 "100011101010",  	 --  2282 	 360 
	 "100011100011",  	 --  2275 	 361 
	 "100011100101",  	 --  2277 	 362 
	 "100011110000",  	 --  2288 	 363 
	 "100100000100",  	 --  2308 	 364 
	 "100100100001",  	 --  2337 	 365 
	 "100101000110",  	 --  2374 	 366 
	 "100101110100",  	 --  2420 	 367 
	 "100110101001",  	 --  2473 	 368 
	 "100111100101",  	 --  2533 	 369 
	 "101000100111",  	 --  2599 	 370 
	 "101001110000",  	 --  2672 	 371 
	 "101010111101",  	 --  2749 	 372 
	 "101100001111",  	 --  2831 	 373 
	 "101101100101",  	 --  2917 	 374 
	 "101110111101",  	 --  3005 	 375 
	 "110000010111",  	 --  3095 	 376 
	 "110001110010",  	 --  3186 	 377 
	 "110011001101",  	 --  3277 	 378 
	 "110100100111",  	 --  3367 	 379 
	 "110101111111",  	 --  3455 	 380 
	 "110111010100",  	 --  3540 	 381 
	 "111000100110",  	 --  3622 	 382 
	 "111001110011",  	 --  3699 	 383 
	 "111010111100",  	 --  3772 	 384 
	 "111011111110",  	 --  3838 	 385 
	 "111100111010",  	 --  3898 	 386 
	 "111101101111",  	 --  3951 	 387 
	 "111110011100",  	 --  3996 	 388 
	 "111111000001",  	 --  4033 	 389 
	 "111111011110",  	 --  4062 	 390 
	 "111111110010",  	 --  4082 	 391 
	 "111111111101",  	 --  4093 	 392 
	 "111111111111",  	 --  4095 	 393 
	 "111111110111",  	 --  4087 	 394 
	 "111111100111",  	 --  4071 	 395 
	 "111111001110",  	 --  4046 	 396 
	 "111110101100",  	 --  4012 	 397 
	 "111110000010",  	 --  3970 	 398 
	 "111101010000",  	 --  3920 	 399 
	 "111100010111",  	 --  3863 	 400 
	 "111011010111",  	 --  3799 	 401 
	 "111010010001",  	 --  3729 	 402 
	 "111001000101",  	 --  3653 	 403 
	 "110111110101",  	 --  3573 	 404 
	 "110110100001",  	 --  3489 	 405 
	 "110101001010",  	 --  3402 	 406 
	 "110011110001",  	 --  3313 	 407 
	 "110010010110",  	 --  3222 	 408 
	 "110000111011",  	 --  3131 	 409 
	 "101111100001",  	 --  3041 	 410 
	 "101110001000",  	 --  2952 	 411 
	 "101100110001",  	 --  2865 	 412 
	 "101011011110",  	 --  2782 	 413 
	 "101010001110",  	 --  2702 	 414 
	 "101001000100",  	 --  2628 	 415 
	 "100111111111",  	 --  2559 	 416 
	 "100111000000",  	 --  2496 	 417 
	 "100110001000",  	 --  2440 	 418 
	 "100101010111",  	 --  2391 	 419 
	 "100100101111",  	 --  2351 	 420 
	 "100100001111",  	 --  2319 	 421 
	 "100011110111",  	 --  2295 	 422 
	 "100011101001",  	 --  2281 	 423 
	 "100011100011",  	 --  2275 	 424 
	 "100011100111",  	 --  2279 	 425 
	 "100011110011",  	 --  2291 	 426 
	 "100100001001",  	 --  2313 	 427 
	 "100100100111",  	 --  2343 	 428 
	 "100101001101",  	 --  2381 	 429 
	 "100101111100",  	 --  2428 	 430 
	 "100110110010",  	 --  2482 	 431 
	 "100111110000",  	 --  2544 	 432 
	 "101000110011",  	 --  2611 	 433 
	 "101001111101",  	 --  2685 	 434 
	 "101011001011",  	 --  2763 	 435 
	 "101100011110",  	 --  2846 	 436 
	 "101101110100",  	 --  2932 	 437 
	 "101111001100",  	 --  3020 	 438 
	 "110000100110",  	 --  3110 	 439 
	 "110010000001",  	 --  3201 	 440 
	 "110011011100",  	 --  3292 	 441 
	 "110100110110",  	 --  3382 	 442 
	 "110110001101",  	 --  3469 	 443 
	 "110111100010",  	 --  3554 	 444 
	 "111000110011",  	 --  3635 	 445 
	 "111010000000",  	 --  3712 	 446 
	 "111011000111",  	 --  3783 	 447 
	 "111100001001",  	 --  3849 	 448 
	 "111101000100",  	 --  3908 	 449 
	 "111101110111",  	 --  3959 	 450 
	 "111110100011",  	 --  4003 	 451 
	 "111111000111",  	 --  4039 	 452 
	 "111111100010",  	 --  4066 	 453 
	 "111111110100",  	 --  4084 	 454 
	 "111111111110",  	 --  4094 	 455 
	 "111111111110",  	 --  4094 	 456 
	 "111111110101",  	 --  4085 	 457 
	 "111111100011",  	 --  4067 	 458 
	 "111111001001",  	 --  4041 	 459 
	 "111110100110",  	 --  4006 	 460 
	 "111101111010",  	 --  3962 	 461 
	 "111101000111",  	 --  3911 	 462 
	 "111100001101",  	 --  3853 	 463 
	 "111011001100",  	 --  3788 	 464 
	 "111010000101",  	 --  3717 	 465 
	 "111000111000",  	 --  3640 	 466 
	 "110111100111",  	 --  3559 	 467 
	 "110110010011",  	 --  3475 	 468 
	 "110100111011",  	 --  3387 	 469 
	 "110011100001",  	 --  3297 	 470 
	 "110010000111",  	 --  3207 	 471 
	 "110000101100",  	 --  3116 	 472 
	 "101111010010",  	 --  3026 	 473 
	 "101101111001",  	 --  2937 	 474 
	 "101100100011",  	 --  2851 	 475 
	 "101011010000",  	 --  2768 	 476 
	 "101010000001",  	 --  2689 	 477 
	 "101000111000",  	 --  2616 	 478 
	 "100111110100",  	 --  2548 	 479 
	 "100110110110",  	 --  2486 	 480 
	 "100101111111",  	 --  2431 	 481 
	 "100101010000",  	 --  2384 	 482 
	 "100100101001",  	 --  2345 	 483 
	 "100100001010",  	 --  2314 	 484 
	 "100011110100",  	 --  2292 	 485 
	 "100011100111",  	 --  2279 	 486 
	 "100011100011",  	 --  2275 	 487 
	 "100011101000",  	 --  2280 	 488 
	 "100011110110",  	 --  2294 	 489 
	 "100100001101",  	 --  2317 	 490 
	 "100100101101",  	 --  2349 	 491 
	 "100101010101",  	 --  2389 	 492 
	 "100110000101",  	 --  2437 	 493 
	 "100110111100",  	 --  2492 	 494 
	 "100111111010",  	 --  2554 	 495 
	 "101000111111",  	 --  2623 	 496 
	 "101010001001",  	 --  2697 	 497 
	 "101011011001",  	 --  2777 	 498 
	 "101100101100",  	 --  2860 	 499 
	 "101110000010",  	 --  2946 	 500 
	 "101111011011",  	 --  3035 	 501 
	 "110000110101",  	 --  3125 	 502 
	 "110010010000",  	 --  3216 	 503 
	 "110011101011",  	 --  3307 	 504 
	 "110101000100",  	 --  3396 	 505 
	 "110110011100",  	 --  3484 	 506 
	 "110111110000",  	 --  3568 	 507 
	 "111001000001",  	 --  3649 	 508 
	 "111010001100",  	 --  3724 	 509 
	 "111011010011",  	 --  3795 	 510 
 	"111100010011");  --  3859 	 511
	begin 
		return tmp;
	end init_rom;
	signal rom : memory_t := init_rom;
begin
	process(clk,ADDR)
		variable addr2 : natural range 0 to 2**m - 1;
	begin
	addr2 := to_integer(unsigned(ADDR));
	if( falling_edge(clk)) then
		q <= rom(addr2);
	end if;
	end process;
end rtl;
