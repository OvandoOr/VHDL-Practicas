library IEEE;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;

entity Comparador_MayorIgual is
	generic(
	n: integer := 8
	);
	port(
	A: 		in std_logic_vector(n-1 downto 0);
	B:		in std_logic_vector(n-1 downto 0);
	MayorIgual:	out std_logic
	);
end Comparador_MayorIgual;

architecture Comparador of Comparador_MayorIgual is
begin
	combinacional: process(A,B)
	begin
		if(A >= B) then
			MayorIgual <= '1';
		else
			MayorIgual <= '0';
		end if;
	end process combinacional;

end Comparador;


















































































































































































































































































































































































































































































































































































