library ieee; 
use ieee.std_logic_1164.all;	
use ieee.numeric_std.all;
entity Rom_Histograma_square is
	generic(
	n: 	integer:= 12;		-- No. de bits informacion
	m:	integer:= 9 		-- No. de bits para datos
	); 
	port 
	(
		CLK		: in std_logic;
		addr	: in std_logic_vector (m-1 downto 0);
		q		: out std_logic_vector((n -1) downto 0)
	);
end Rom_Histograma_square;
architecture rtl of Rom_Histograma_square is
	subtype word_t is std_logic_vector((n-1) downto 0);
	type memory_t is array(0 to (2**m)-1 ) of word_t;
	function init_rom
		return memory_t is 
		variable tmp : memory_t :=(
	 "111111111111",  	 --  4095 	 0 
	 "111111111111",  	 --  4095 	 1 
	 "111111111111",  	 --  4095 	 2 
	 "111111111111",  	 --  4095 	 3 
	 "111111111111",  	 --  4095 	 4 
	 "111111111111",  	 --  4095 	 5 
	 "111111111111",  	 --  4095 	 6 
	 "111111111111",  	 --  4095 	 7 
	 "111111111111",  	 --  4095 	 8 
	 "111111111111",  	 --  4095 	 9 
	 "111111111111",  	 --  4095 	 10 
	 "111111111111",  	 --  4095 	 11 
	 "111111111111",  	 --  4095 	 12 
	 "111111111111",  	 --  4095 	 13 
	 "111111111111",  	 --  4095 	 14 
	 "111111111111",  	 --  4095 	 15 
	 "111111111111",  	 --  4095 	 16 
	 "111111111111",  	 --  4095 	 17 
	 "111111111111",  	 --  4095 	 18 
	 "111111111111",  	 --  4095 	 19 
	 "111111111111",  	 --  4095 	 20 
	 "111111111111",  	 --  4095 	 21 
	 "111111111111",  	 --  4095 	 22 
	 "111111111111",  	 --  4095 	 23 
	 "111111111111",  	 --  4095 	 24 
	 "111111111111",  	 --  4095 	 25 
	 "111111111111",  	 --  4095 	 26 
	 "111111111111",  	 --  4095 	 27 
	 "111111111111",  	 --  4095 	 28 
	 "111111111111",  	 --  4095 	 29 
	 "111111111111",  	 --  4095 	 30 
	 "111111111111",  	 --  4095 	 31 
	 "100011100011",  	 --  2275 	 32 
	 "100011100011",  	 --  2275 	 33 
	 "100011100011",  	 --  2275 	 34 
	 "100011100011",  	 --  2275 	 35 
	 "100011100011",  	 --  2275 	 36 
	 "100011100011",  	 --  2275 	 37 
	 "100011100011",  	 --  2275 	 38 
	 "100011100011",  	 --  2275 	 39 
	 "100011100011",  	 --  2275 	 40 
	 "100011100011",  	 --  2275 	 41 
	 "100011100011",  	 --  2275 	 42 
	 "100011100011",  	 --  2275 	 43 
	 "100011100011",  	 --  2275 	 44 
	 "100011100011",  	 --  2275 	 45 
	 "100011100011",  	 --  2275 	 46 
	 "100011100011",  	 --  2275 	 47 
	 "100011100011",  	 --  2275 	 48 
	 "100011100011",  	 --  2275 	 49 
	 "100011100011",  	 --  2275 	 50 
	 "100011100011",  	 --  2275 	 51 
	 "100011100011",  	 --  2275 	 52 
	 "100011100011",  	 --  2275 	 53 
	 "100011100011",  	 --  2275 	 54 
	 "100011100011",  	 --  2275 	 55 
	 "100011100011",  	 --  2275 	 56 
	 "100011100011",  	 --  2275 	 57 
	 "100011100011",  	 --  2275 	 58 
	 "100011100011",  	 --  2275 	 59 
	 "100011100011",  	 --  2275 	 60 
	 "100011100011",  	 --  2275 	 61 
	 "100011100011",  	 --  2275 	 62 
	 "111111111111",  	 --  4095 	 63 
	 "111111111111",  	 --  4095 	 64 
	 "111111111111",  	 --  4095 	 65 
	 "111111111111",  	 --  4095 	 66 
	 "111111111111",  	 --  4095 	 67 
	 "111111111111",  	 --  4095 	 68 
	 "111111111111",  	 --  4095 	 69 
	 "111111111111",  	 --  4095 	 70 
	 "111111111111",  	 --  4095 	 71 
	 "111111111111",  	 --  4095 	 72 
	 "111111111111",  	 --  4095 	 73 
	 "111111111111",  	 --  4095 	 74 
	 "111111111111",  	 --  4095 	 75 
	 "111111111111",  	 --  4095 	 76 
	 "111111111111",  	 --  4095 	 77 
	 "111111111111",  	 --  4095 	 78 
	 "111111111111",  	 --  4095 	 79 
	 "111111111111",  	 --  4095 	 80 
	 "111111111111",  	 --  4095 	 81 
	 "111111111111",  	 --  4095 	 82 
	 "111111111111",  	 --  4095 	 83 
	 "111111111111",  	 --  4095 	 84 
	 "111111111111",  	 --  4095 	 85 
	 "111111111111",  	 --  4095 	 86 
	 "111111111111",  	 --  4095 	 87 
	 "111111111111",  	 --  4095 	 88 
	 "111111111111",  	 --  4095 	 89 
	 "111111111111",  	 --  4095 	 90 
	 "111111111111",  	 --  4095 	 91 
	 "111111111111",  	 --  4095 	 92 
	 "111111111111",  	 --  4095 	 93 
	 "111111111111",  	 --  4095 	 94 
	 "100011100011",  	 --  2275 	 95 
	 "100011100011",  	 --  2275 	 96 
	 "100011100011",  	 --  2275 	 97 
	 "100011100011",  	 --  2275 	 98 
	 "100011100011",  	 --  2275 	 99 
	 "100011100011",  	 --  2275 	 100 
	 "100011100011",  	 --  2275 	 101 
	 "100011100011",  	 --  2275 	 102 
	 "100011100011",  	 --  2275 	 103 
	 "100011100011",  	 --  2275 	 104 
	 "100011100011",  	 --  2275 	 105 
	 "100011100011",  	 --  2275 	 106 
	 "100011100011",  	 --  2275 	 107 
	 "100011100011",  	 --  2275 	 108 
	 "100011100011",  	 --  2275 	 109 
	 "100011100011",  	 --  2275 	 110 
	 "100011100011",  	 --  2275 	 111 
	 "100011100011",  	 --  2275 	 112 
	 "100011100011",  	 --  2275 	 113 
	 "100011100011",  	 --  2275 	 114 
	 "100011100011",  	 --  2275 	 115 
	 "100011100011",  	 --  2275 	 116 
	 "100011100011",  	 --  2275 	 117 
	 "100011100011",  	 --  2275 	 118 
	 "100011100011",  	 --  2275 	 119 
	 "100011100011",  	 --  2275 	 120 
	 "100011100011",  	 --  2275 	 121 
	 "100011100011",  	 --  2275 	 122 
	 "100011100011",  	 --  2275 	 123 
	 "100011100011",  	 --  2275 	 124 
	 "100011100011",  	 --  2275 	 125 
	 "111111111111",  	 --  4095 	 126 
	 "111111111111",  	 --  4095 	 127 
	 "111111111111",  	 --  4095 	 128 
	 "111111111111",  	 --  4095 	 129 
	 "111111111111",  	 --  4095 	 130 
	 "111111111111",  	 --  4095 	 131 
	 "111111111111",  	 --  4095 	 132 
	 "111111111111",  	 --  4095 	 133 
	 "111111111111",  	 --  4095 	 134 
	 "111111111111",  	 --  4095 	 135 
	 "111111111111",  	 --  4095 	 136 
	 "111111111111",  	 --  4095 	 137 
	 "111111111111",  	 --  4095 	 138 
	 "111111111111",  	 --  4095 	 139 
	 "111111111111",  	 --  4095 	 140 
	 "111111111111",  	 --  4095 	 141 
	 "111111111111",  	 --  4095 	 142 
	 "111111111111",  	 --  4095 	 143 
	 "111111111111",  	 --  4095 	 144 
	 "111111111111",  	 --  4095 	 145 
	 "111111111111",  	 --  4095 	 146 
	 "111111111111",  	 --  4095 	 147 
	 "111111111111",  	 --  4095 	 148 
	 "111111111111",  	 --  4095 	 149 
	 "111111111111",  	 --  4095 	 150 
	 "111111111111",  	 --  4095 	 151 
	 "111111111111",  	 --  4095 	 152 
	 "111111111111",  	 --  4095 	 153 
	 "111111111111",  	 --  4095 	 154 
	 "111111111111",  	 --  4095 	 155 
	 "111111111111",  	 --  4095 	 156 
	 "111111111111",  	 --  4095 	 157 
	 "100011100011",  	 --  2275 	 158 
	 "100011100011",  	 --  2275 	 159 
	 "100011100011",  	 --  2275 	 160 
	 "100011100011",  	 --  2275 	 161 
	 "100011100011",  	 --  2275 	 162 
	 "100011100011",  	 --  2275 	 163 
	 "100011100011",  	 --  2275 	 164 
	 "100011100011",  	 --  2275 	 165 
	 "100011100011",  	 --  2275 	 166 
	 "100011100011",  	 --  2275 	 167 
	 "100011100011",  	 --  2275 	 168 
	 "100011100011",  	 --  2275 	 169 
	 "100011100011",  	 --  2275 	 170 
	 "100011100011",  	 --  2275 	 171 
	 "100011100011",  	 --  2275 	 172 
	 "100011100011",  	 --  2275 	 173 
	 "100011100011",  	 --  2275 	 174 
	 "100011100011",  	 --  2275 	 175 
	 "100011100011",  	 --  2275 	 176 
	 "100011100011",  	 --  2275 	 177 
	 "100011100011",  	 --  2275 	 178 
	 "100011100011",  	 --  2275 	 179 
	 "100011100011",  	 --  2275 	 180 
	 "100011100011",  	 --  2275 	 181 
	 "100011100011",  	 --  2275 	 182 
	 "100011100011",  	 --  2275 	 183 
	 "100011100011",  	 --  2275 	 184 
	 "100011100011",  	 --  2275 	 185 
	 "100011100011",  	 --  2275 	 186 
	 "100011100011",  	 --  2275 	 187 
	 "100011100011",  	 --  2275 	 188 
	 "111111111111",  	 --  4095 	 189 
	 "111111111111",  	 --  4095 	 190 
	 "111111111111",  	 --  4095 	 191 
	 "111111111111",  	 --  4095 	 192 
	 "111111111111",  	 --  4095 	 193 
	 "111111111111",  	 --  4095 	 194 
	 "111111111111",  	 --  4095 	 195 
	 "111111111111",  	 --  4095 	 196 
	 "111111111111",  	 --  4095 	 197 
	 "111111111111",  	 --  4095 	 198 
	 "111111111111",  	 --  4095 	 199 
	 "111111111111",  	 --  4095 	 200 
	 "111111111111",  	 --  4095 	 201 
	 "111111111111",  	 --  4095 	 202 
	 "111111111111",  	 --  4095 	 203 
	 "111111111111",  	 --  4095 	 204 
	 "111111111111",  	 --  4095 	 205 
	 "111111111111",  	 --  4095 	 206 
	 "111111111111",  	 --  4095 	 207 
	 "111111111111",  	 --  4095 	 208 
	 "111111111111",  	 --  4095 	 209 
	 "111111111111",  	 --  4095 	 210 
	 "111111111111",  	 --  4095 	 211 
	 "111111111111",  	 --  4095 	 212 
	 "111111111111",  	 --  4095 	 213 
	 "111111111111",  	 --  4095 	 214 
	 "111111111111",  	 --  4095 	 215 
	 "111111111111",  	 --  4095 	 216 
	 "111111111111",  	 --  4095 	 217 
	 "111111111111",  	 --  4095 	 218 
	 "111111111111",  	 --  4095 	 219 
	 "100011100011",  	 --  2275 	 220 
	 "100011100011",  	 --  2275 	 221 
	 "100011100011",  	 --  2275 	 222 
	 "100011100011",  	 --  2275 	 223 
	 "100011100011",  	 --  2275 	 224 
	 "100011100011",  	 --  2275 	 225 
	 "100011100011",  	 --  2275 	 226 
	 "100011100011",  	 --  2275 	 227 
	 "100011100011",  	 --  2275 	 228 
	 "100011100011",  	 --  2275 	 229 
	 "100011100011",  	 --  2275 	 230 
	 "100011100011",  	 --  2275 	 231 
	 "100011100011",  	 --  2275 	 232 
	 "100011100011",  	 --  2275 	 233 
	 "100011100011",  	 --  2275 	 234 
	 "100011100011",  	 --  2275 	 235 
	 "100011100011",  	 --  2275 	 236 
	 "100011100011",  	 --  2275 	 237 
	 "100011100011",  	 --  2275 	 238 
	 "100011100011",  	 --  2275 	 239 
	 "100011100011",  	 --  2275 	 240 
	 "100011100011",  	 --  2275 	 241 
	 "100011100011",  	 --  2275 	 242 
	 "100011100011",  	 --  2275 	 243 
	 "100011100011",  	 --  2275 	 244 
	 "100011100011",  	 --  2275 	 245 
	 "100011100011",  	 --  2275 	 246 
	 "100011100011",  	 --  2275 	 247 
	 "100011100011",  	 --  2275 	 248 
	 "100011100011",  	 --  2275 	 249 
	 "100011100011",  	 --  2275 	 250 
	 "100011100011",  	 --  2275 	 251 
	 "111111111111",  	 --  4095 	 252 
	 "111111111111",  	 --  4095 	 253 
	 "111111111111",  	 --  4095 	 254 
	 "111111111111",  	 --  4095 	 255 
	 "111111111111",  	 --  4095 	 256 
	 "111111111111",  	 --  4095 	 257 
	 "111111111111",  	 --  4095 	 258 
	 "111111111111",  	 --  4095 	 259 
	 "111111111111",  	 --  4095 	 260 
	 "111111111111",  	 --  4095 	 261 
	 "111111111111",  	 --  4095 	 262 
	 "111111111111",  	 --  4095 	 263 
	 "111111111111",  	 --  4095 	 264 
	 "111111111111",  	 --  4095 	 265 
	 "111111111111",  	 --  4095 	 266 
	 "111111111111",  	 --  4095 	 267 
	 "111111111111",  	 --  4095 	 268 
	 "111111111111",  	 --  4095 	 269 
	 "111111111111",  	 --  4095 	 270 
	 "111111111111",  	 --  4095 	 271 
	 "111111111111",  	 --  4095 	 272 
	 "111111111111",  	 --  4095 	 273 
	 "111111111111",  	 --  4095 	 274 
	 "111111111111",  	 --  4095 	 275 
	 "111111111111",  	 --  4095 	 276 
	 "111111111111",  	 --  4095 	 277 
	 "111111111111",  	 --  4095 	 278 
	 "111111111111",  	 --  4095 	 279 
	 "111111111111",  	 --  4095 	 280 
	 "111111111111",  	 --  4095 	 281 
	 "111111111111",  	 --  4095 	 282 
	 "100011100011",  	 --  2275 	 283 
	 "100011100011",  	 --  2275 	 284 
	 "100011100011",  	 --  2275 	 285 
	 "100011100011",  	 --  2275 	 286 
	 "100011100011",  	 --  2275 	 287 
	 "100011100011",  	 --  2275 	 288 
	 "100011100011",  	 --  2275 	 289 
	 "100011100011",  	 --  2275 	 290 
	 "100011100011",  	 --  2275 	 291 
	 "100011100011",  	 --  2275 	 292 
	 "100011100011",  	 --  2275 	 293 
	 "100011100011",  	 --  2275 	 294 
	 "100011100011",  	 --  2275 	 295 
	 "100011100011",  	 --  2275 	 296 
	 "100011100011",  	 --  2275 	 297 
	 "100011100011",  	 --  2275 	 298 
	 "100011100011",  	 --  2275 	 299 
	 "100011100011",  	 --  2275 	 300 
	 "100011100011",  	 --  2275 	 301 
	 "100011100011",  	 --  2275 	 302 
	 "100011100011",  	 --  2275 	 303 
	 "100011100011",  	 --  2275 	 304 
	 "100011100011",  	 --  2275 	 305 
	 "100011100011",  	 --  2275 	 306 
	 "100011100011",  	 --  2275 	 307 
	 "100011100011",  	 --  2275 	 308 
	 "100011100011",  	 --  2275 	 309 
	 "100011100011",  	 --  2275 	 310 
	 "100011100011",  	 --  2275 	 311 
	 "100011100011",  	 --  2275 	 312 
	 "100011100011",  	 --  2275 	 313 
	 "100011100011",  	 --  2275 	 314 
	 "111111111111",  	 --  4095 	 315 
	 "111111111111",  	 --  4095 	 316 
	 "111111111111",  	 --  4095 	 317 
	 "111111111111",  	 --  4095 	 318 
	 "111111111111",  	 --  4095 	 319 
	 "111111111111",  	 --  4095 	 320 
	 "111111111111",  	 --  4095 	 321 
	 "111111111111",  	 --  4095 	 322 
	 "111111111111",  	 --  4095 	 323 
	 "111111111111",  	 --  4095 	 324 
	 "111111111111",  	 --  4095 	 325 
	 "111111111111",  	 --  4095 	 326 
	 "111111111111",  	 --  4095 	 327 
	 "111111111111",  	 --  4095 	 328 
	 "111111111111",  	 --  4095 	 329 
	 "111111111111",  	 --  4095 	 330 
	 "111111111111",  	 --  4095 	 331 
	 "111111111111",  	 --  4095 	 332 
	 "111111111111",  	 --  4095 	 333 
	 "111111111111",  	 --  4095 	 334 
	 "111111111111",  	 --  4095 	 335 
	 "111111111111",  	 --  4095 	 336 
	 "111111111111",  	 --  4095 	 337 
	 "111111111111",  	 --  4095 	 338 
	 "111111111111",  	 --  4095 	 339 
	 "111111111111",  	 --  4095 	 340 
	 "111111111111",  	 --  4095 	 341 
	 "111111111111",  	 --  4095 	 342 
	 "111111111111",  	 --  4095 	 343 
	 "111111111111",  	 --  4095 	 344 
	 "111111111111",  	 --  4095 	 345 
	 "100011100011",  	 --  2275 	 346 
	 "100011100011",  	 --  2275 	 347 
	 "100011100011",  	 --  2275 	 348 
	 "100011100011",  	 --  2275 	 349 
	 "100011100011",  	 --  2275 	 350 
	 "100011100011",  	 --  2275 	 351 
	 "100011100011",  	 --  2275 	 352 
	 "100011100011",  	 --  2275 	 353 
	 "100011100011",  	 --  2275 	 354 
	 "100011100011",  	 --  2275 	 355 
	 "100011100011",  	 --  2275 	 356 
	 "100011100011",  	 --  2275 	 357 
	 "100011100011",  	 --  2275 	 358 
	 "100011100011",  	 --  2275 	 359 
	 "100011100011",  	 --  2275 	 360 
	 "100011100011",  	 --  2275 	 361 
	 "100011100011",  	 --  2275 	 362 
	 "100011100011",  	 --  2275 	 363 
	 "100011100011",  	 --  2275 	 364 
	 "100011100011",  	 --  2275 	 365 
	 "100011100011",  	 --  2275 	 366 
	 "100011100011",  	 --  2275 	 367 
	 "100011100011",  	 --  2275 	 368 
	 "100011100011",  	 --  2275 	 369 
	 "100011100011",  	 --  2275 	 370 
	 "100011100011",  	 --  2275 	 371 
	 "100011100011",  	 --  2275 	 372 
	 "100011100011",  	 --  2275 	 373 
	 "100011100011",  	 --  2275 	 374 
	 "100011100011",  	 --  2275 	 375 
	 "100011100011",  	 --  2275 	 376 
	 "111111111111",  	 --  4095 	 377 
	 "111111111111",  	 --  4095 	 378 
	 "111111111111",  	 --  4095 	 379 
	 "111111111111",  	 --  4095 	 380 
	 "111111111111",  	 --  4095 	 381 
	 "111111111111",  	 --  4095 	 382 
	 "111111111111",  	 --  4095 	 383 
	 "111111111111",  	 --  4095 	 384 
	 "111111111111",  	 --  4095 	 385 
	 "111111111111",  	 --  4095 	 386 
	 "111111111111",  	 --  4095 	 387 
	 "111111111111",  	 --  4095 	 388 
	 "111111111111",  	 --  4095 	 389 
	 "111111111111",  	 --  4095 	 390 
	 "111111111111",  	 --  4095 	 391 
	 "111111111111",  	 --  4095 	 392 
	 "111111111111",  	 --  4095 	 393 
	 "111111111111",  	 --  4095 	 394 
	 "111111111111",  	 --  4095 	 395 
	 "111111111111",  	 --  4095 	 396 
	 "111111111111",  	 --  4095 	 397 
	 "111111111111",  	 --  4095 	 398 
	 "111111111111",  	 --  4095 	 399 
	 "111111111111",  	 --  4095 	 400 
	 "111111111111",  	 --  4095 	 401 
	 "111111111111",  	 --  4095 	 402 
	 "111111111111",  	 --  4095 	 403 
	 "111111111111",  	 --  4095 	 404 
	 "111111111111",  	 --  4095 	 405 
	 "111111111111",  	 --  4095 	 406 
	 "111111111111",  	 --  4095 	 407 
	 "111111111111",  	 --  4095 	 408 
	 "100011100011",  	 --  2275 	 409 
	 "100011100011",  	 --  2275 	 410 
	 "100011100011",  	 --  2275 	 411 
	 "100011100011",  	 --  2275 	 412 
	 "100011100011",  	 --  2275 	 413 
	 "100011100011",  	 --  2275 	 414 
	 "100011100011",  	 --  2275 	 415 
	 "100011100011",  	 --  2275 	 416 
	 "100011100011",  	 --  2275 	 417 
	 "100011100011",  	 --  2275 	 418 
	 "100011100011",  	 --  2275 	 419 
	 "100011100011",  	 --  2275 	 420 
	 "100011100011",  	 --  2275 	 421 
	 "100011100011",  	 --  2275 	 422 
	 "100011100011",  	 --  2275 	 423 
	 "100011100011",  	 --  2275 	 424 
	 "100011100011",  	 --  2275 	 425 
	 "100011100011",  	 --  2275 	 426 
	 "100011100011",  	 --  2275 	 427 
	 "100011100011",  	 --  2275 	 428 
	 "100011100011",  	 --  2275 	 429 
	 "100011100011",  	 --  2275 	 430 
	 "100011100011",  	 --  2275 	 431 
	 "100011100011",  	 --  2275 	 432 
	 "100011100011",  	 --  2275 	 433 
	 "100011100011",  	 --  2275 	 434 
	 "100011100011",  	 --  2275 	 435 
	 "100011100011",  	 --  2275 	 436 
	 "100011100011",  	 --  2275 	 437 
	 "100011100011",  	 --  2275 	 438 
	 "100011100011",  	 --  2275 	 439 
	 "111111111111",  	 --  4095 	 440 
	 "111111111111",  	 --  4095 	 441 
	 "111111111111",  	 --  4095 	 442 
	 "111111111111",  	 --  4095 	 443 
	 "111111111111",  	 --  4095 	 444 
	 "111111111111",  	 --  4095 	 445 
	 "111111111111",  	 --  4095 	 446 
	 "111111111111",  	 --  4095 	 447 
	 "111111111111",  	 --  4095 	 448 
	 "111111111111",  	 --  4095 	 449 
	 "111111111111",  	 --  4095 	 450 
	 "111111111111",  	 --  4095 	 451 
	 "111111111111",  	 --  4095 	 452 
	 "111111111111",  	 --  4095 	 453 
	 "111111111111",  	 --  4095 	 454 
	 "111111111111",  	 --  4095 	 455 
	 "111111111111",  	 --  4095 	 456 
	 "111111111111",  	 --  4095 	 457 
	 "111111111111",  	 --  4095 	 458 
	 "111111111111",  	 --  4095 	 459 
	 "111111111111",  	 --  4095 	 460 
	 "111111111111",  	 --  4095 	 461 
	 "111111111111",  	 --  4095 	 462 
	 "111111111111",  	 --  4095 	 463 
	 "111111111111",  	 --  4095 	 464 
	 "111111111111",  	 --  4095 	 465 
	 "111111111111",  	 --  4095 	 466 
	 "111111111111",  	 --  4095 	 467 
	 "111111111111",  	 --  4095 	 468 
	 "111111111111",  	 --  4095 	 469 
	 "111111111111",  	 --  4095 	 470 
	 "111111111111",  	 --  4095 	 471 
	 "100011100011",  	 --  2275 	 472 
	 "100011100011",  	 --  2275 	 473 
	 "100011100011",  	 --  2275 	 474 
	 "100011100011",  	 --  2275 	 475 
	 "100011100011",  	 --  2275 	 476 
	 "100011100011",  	 --  2275 	 477 
	 "100011100011",  	 --  2275 	 478 
	 "100011100011",  	 --  2275 	 479 
	 "100011100011",  	 --  2275 	 480 
	 "100011100011",  	 --  2275 	 481 
	 "100011100011",  	 --  2275 	 482 
	 "100011100011",  	 --  2275 	 483 
	 "100011100011",  	 --  2275 	 484 
	 "100011100011",  	 --  2275 	 485 
	 "100011100011",  	 --  2275 	 486 
	 "100011100011",  	 --  2275 	 487 
	 "100011100011",  	 --  2275 	 488 
	 "100011100011",  	 --  2275 	 489 
	 "100011100011",  	 --  2275 	 490 
	 "100011100011",  	 --  2275 	 491 
	 "100011100011",  	 --  2275 	 492 
	 "100011100011",  	 --  2275 	 493 
	 "100011100011",  	 --  2275 	 494 
	 "100011100011",  	 --  2275 	 495 
	 "100011100011",  	 --  2275 	 496 
	 "100011100011",  	 --  2275 	 497 
	 "100011100011",  	 --  2275 	 498 
	 "100011100011",  	 --  2275 	 499 
	 "100011100011",  	 --  2275 	 500 
	 "100011100011",  	 --  2275 	 501 
	 "100011100011",  	 --  2275 	 502 
	 "111111111111",  	 --  4095 	 503 
	 "111111111111",  	 --  4095 	 504 
	 "111111111111",  	 --  4095 	 505 
	 "111111111111",  	 --  4095 	 506 
	 "111111111111",  	 --  4095 	 507 
	 "111111111111",  	 --  4095 	 508 
	 "111111111111",  	 --  4095 	 509 
	 "111111111111",  	 --  4095 	 510 
 	"111111111111");  --  4095 	 511
	begin 
		return tmp;
	end init_rom;
	signal rom : memory_t := init_rom;
begin
	process(clk,ADDR)
		variable addr2 : natural range 0 to 2**m - 1;
	begin
	addr2 := to_integer(unsigned(ADDR));
	if( falling_edge(clk)) then
		q <= rom(addr2);
	end if;
	end process;
end rtl;
