library ieee; 
use ieee.std_logic_1164.all;	
use ieee.numeric_std.all;
entity Rom_Histograma_sawtooth is
	generic(
	n: 	integer:= 12;		-- No. de bits informacion
	m:	integer:= 9 		-- No. de bits para datos
	); 
	port 
	(
		CLK		: in std_logic;
		addr	: in std_logic_vector (m-1 downto 0);
		q		: out std_logic_vector((n -1) downto 0)
	);
end Rom_Histograma_sawtooth;
architecture rtl of Rom_Histograma_sawtooth is
	subtype word_t is std_logic_vector((n-1) downto 0);
	type memory_t is array(0 to (2**m)-1 ) of word_t;
	function init_rom
		return memory_t is 
		variable tmp : memory_t :=(
	 "100011100011",  	 --  2275 	 0 
	 "100100000000",  	 --  2304 	 1 
	 "100100011101",  	 --  2333 	 2 
	 "100100111010",  	 --  2362 	 3 
	 "100101010111",  	 --  2391 	 4 
	 "100101110100",  	 --  2420 	 5 
	 "100110010001",  	 --  2449 	 6 
	 "100110101110",  	 --  2478 	 7 
	 "100111001011",  	 --  2507 	 8 
	 "100111101000",  	 --  2536 	 9 
	 "101000000101",  	 --  2565 	 10 
	 "101000100010",  	 --  2594 	 11 
	 "101000111111",  	 --  2623 	 12 
	 "101001011100",  	 --  2652 	 13 
	 "101001111001",  	 --  2681 	 14 
	 "101010010101",  	 --  2709 	 15 
	 "101010110010",  	 --  2738 	 16 
	 "101011001111",  	 --  2767 	 17 
	 "101011101100",  	 --  2796 	 18 
	 "101100001001",  	 --  2825 	 19 
	 "101100100110",  	 --  2854 	 20 
	 "101101000011",  	 --  2883 	 21 
	 "101101100000",  	 --  2912 	 22 
	 "101101111101",  	 --  2941 	 23 
	 "101110011010",  	 --  2970 	 24 
	 "101110110111",  	 --  2999 	 25 
	 "101111010100",  	 --  3028 	 26 
	 "101111110001",  	 --  3057 	 27 
	 "110000001110",  	 --  3086 	 28 
	 "110000101011",  	 --  3115 	 29 
	 "110001001000",  	 --  3144 	 30 
	 "110001100101",  	 --  3173 	 31 
	 "110010000010",  	 --  3202 	 32 
	 "110010011111",  	 --  3231 	 33 
	 "110010111100",  	 --  3260 	 34 
	 "110011011001",  	 --  3289 	 35 
	 "110011110110",  	 --  3318 	 36 
	 "110100010011",  	 --  3347 	 37 
	 "110100110000",  	 --  3376 	 38 
	 "110101001101",  	 --  3405 	 39 
	 "110101101010",  	 --  3434 	 40 
	 "110110000111",  	 --  3463 	 41 
	 "110110100100",  	 --  3492 	 42 
	 "110111000001",  	 --  3521 	 43 
	 "110111011110",  	 --  3550 	 44 
	 "110111111010",  	 --  3578 	 45 
	 "111000010111",  	 --  3607 	 46 
	 "111000110100",  	 --  3636 	 47 
	 "111001010001",  	 --  3665 	 48 
	 "111001101110",  	 --  3694 	 49 
	 "111010001011",  	 --  3723 	 50 
	 "111010101000",  	 --  3752 	 51 
	 "111011000101",  	 --  3781 	 52 
	 "111011100010",  	 --  3810 	 53 
	 "111011111111",  	 --  3839 	 54 
	 "111100011100",  	 --  3868 	 55 
	 "111100111001",  	 --  3897 	 56 
	 "111101010110",  	 --  3926 	 57 
	 "111101110011",  	 --  3955 	 58 
	 "111110010000",  	 --  3984 	 59 
	 "111110101101",  	 --  4013 	 60 
	 "111111001010",  	 --  4042 	 61 
	 "111111100111",  	 --  4071 	 62 
	 "100011101000",  	 --  2280 	 63 
	 "100100000101",  	 --  2309 	 64 
	 "100100100010",  	 --  2338 	 65 
	 "100100111111",  	 --  2367 	 66 
	 "100101011100",  	 --  2396 	 67 
	 "100101111001",  	 --  2425 	 68 
	 "100110010110",  	 --  2454 	 69 
	 "100110110011",  	 --  2483 	 70 
	 "100111010000",  	 --  2512 	 71 
	 "100111101101",  	 --  2541 	 72 
	 "101000001010",  	 --  2570 	 73 
	 "101000100110",  	 --  2598 	 74 
	 "101001000011",  	 --  2627 	 75 
	 "101001100000",  	 --  2656 	 76 
	 "101001111101",  	 --  2685 	 77 
	 "101010011010",  	 --  2714 	 78 
	 "101010110111",  	 --  2743 	 79 
	 "101011010100",  	 --  2772 	 80 
	 "101011110001",  	 --  2801 	 81 
	 "101100001110",  	 --  2830 	 82 
	 "101100101011",  	 --  2859 	 83 
	 "101101001000",  	 --  2888 	 84 
	 "101101100101",  	 --  2917 	 85 
	 "101110000010",  	 --  2946 	 86 
	 "101110011111",  	 --  2975 	 87 
	 "101110111100",  	 --  3004 	 88 
	 "101111011001",  	 --  3033 	 89 
	 "101111110110",  	 --  3062 	 90 
	 "110000010011",  	 --  3091 	 91 
	 "110000110000",  	 --  3120 	 92 
	 "110001001101",  	 --  3149 	 93 
	 "110001101010",  	 --  3178 	 94 
	 "110010000111",  	 --  3207 	 95 
	 "110010100100",  	 --  3236 	 96 
	 "110011000001",  	 --  3265 	 97 
	 "110011011110",  	 --  3294 	 98 
	 "110011111011",  	 --  3323 	 99 
	 "110100011000",  	 --  3352 	 100 
	 "110100110101",  	 --  3381 	 101 
	 "110101010010",  	 --  3410 	 102 
	 "110101101111",  	 --  3439 	 103 
	 "110110001011",  	 --  3467 	 104 
	 "110110101000",  	 --  3496 	 105 
	 "110111000101",  	 --  3525 	 106 
	 "110111100010",  	 --  3554 	 107 
	 "110111111111",  	 --  3583 	 108 
	 "111000011100",  	 --  3612 	 109 
	 "111000111001",  	 --  3641 	 110 
	 "111001010110",  	 --  3670 	 111 
	 "111001110011",  	 --  3699 	 112 
	 "111010010000",  	 --  3728 	 113 
	 "111010101101",  	 --  3757 	 114 
	 "111011001010",  	 --  3786 	 115 
	 "111011100111",  	 --  3815 	 116 
	 "111100000100",  	 --  3844 	 117 
	 "111100100001",  	 --  3873 	 118 
	 "111100111110",  	 --  3902 	 119 
	 "111101011011",  	 --  3931 	 120 
	 "111101111000",  	 --  3960 	 121 
	 "111110010101",  	 --  3989 	 122 
	 "111110110010",  	 --  4018 	 123 
	 "111111001111",  	 --  4047 	 124 
	 "111111101100",  	 --  4076 	 125 
	 "100011101101",  	 --  2285 	 126 
	 "100100001010",  	 --  2314 	 127 
	 "100100100111",  	 --  2343 	 128 
	 "100101000100",  	 --  2372 	 129 
	 "100101100001",  	 --  2401 	 130 
	 "100101111110",  	 --  2430 	 131 
	 "100110011011",  	 --  2459 	 132 
	 "100110111000",  	 --  2488 	 133 
	 "100111010100",  	 --  2516 	 134 
	 "100111110001",  	 --  2545 	 135 
	 "101000001110",  	 --  2574 	 136 
	 "101000101011",  	 --  2603 	 137 
	 "101001001000",  	 --  2632 	 138 
	 "101001100101",  	 --  2661 	 139 
	 "101010000010",  	 --  2690 	 140 
	 "101010011111",  	 --  2719 	 141 
	 "101010111100",  	 --  2748 	 142 
	 "101011011001",  	 --  2777 	 143 
	 "101011110110",  	 --  2806 	 144 
	 "101100010011",  	 --  2835 	 145 
	 "101100110000",  	 --  2864 	 146 
	 "101101001101",  	 --  2893 	 147 
	 "101101101010",  	 --  2922 	 148 
	 "101110000111",  	 --  2951 	 149 
	 "101110100100",  	 --  2980 	 150 
	 "101111000001",  	 --  3009 	 151 
	 "101111011110",  	 --  3038 	 152 
	 "101111111011",  	 --  3067 	 153 
	 "110000011000",  	 --  3096 	 154 
	 "110000110101",  	 --  3125 	 155 
	 "110001010010",  	 --  3154 	 156 
	 "110001101111",  	 --  3183 	 157 
	 "110010001100",  	 --  3212 	 158 
	 "110010101001",  	 --  3241 	 159 
	 "110011000110",  	 --  3270 	 160 
	 "110011100011",  	 --  3299 	 161 
	 "110100000000",  	 --  3328 	 162 
	 "110100011100",  	 --  3356 	 163 
	 "110100111001",  	 --  3385 	 164 
	 "110101010110",  	 --  3414 	 165 
	 "110101110011",  	 --  3443 	 166 
	 "110110010000",  	 --  3472 	 167 
	 "110110101101",  	 --  3501 	 168 
	 "110111001010",  	 --  3530 	 169 
	 "110111100111",  	 --  3559 	 170 
	 "111000000100",  	 --  3588 	 171 
	 "111000100001",  	 --  3617 	 172 
	 "111000111110",  	 --  3646 	 173 
	 "111001011011",  	 --  3675 	 174 
	 "111001111000",  	 --  3704 	 175 
	 "111010010101",  	 --  3733 	 176 
	 "111010110010",  	 --  3762 	 177 
	 "111011001111",  	 --  3791 	 178 
	 "111011101100",  	 --  3820 	 179 
	 "111100001001",  	 --  3849 	 180 
	 "111100100110",  	 --  3878 	 181 
	 "111101000011",  	 --  3907 	 182 
	 "111101100000",  	 --  3936 	 183 
	 "111101111101",  	 --  3965 	 184 
	 "111110011010",  	 --  3994 	 185 
	 "111110110111",  	 --  4023 	 186 
	 "111111010100",  	 --  4052 	 187 
	 "111111110001",  	 --  4081 	 188 
	 "100011110010",  	 --  2290 	 189 
	 "100100001111",  	 --  2319 	 190 
	 "100100101100",  	 --  2348 	 191 
	 "100101001001",  	 --  2377 	 192 
	 "100101100101",  	 --  2405 	 193 
	 "100110000010",  	 --  2434 	 194 
	 "100110011111",  	 --  2463 	 195 
	 "100110111100",  	 --  2492 	 196 
	 "100111011001",  	 --  2521 	 197 
	 "100111110110",  	 --  2550 	 198 
	 "101000010011",  	 --  2579 	 199 
	 "101000110000",  	 --  2608 	 200 
	 "101001001101",  	 --  2637 	 201 
	 "101001101010",  	 --  2666 	 202 
	 "101010000111",  	 --  2695 	 203 
	 "101010100100",  	 --  2724 	 204 
	 "101011000001",  	 --  2753 	 205 
	 "101011011110",  	 --  2782 	 206 
	 "101011111011",  	 --  2811 	 207 
	 "101100011000",  	 --  2840 	 208 
	 "101100110101",  	 --  2869 	 209 
	 "101101010010",  	 --  2898 	 210 
	 "101101101111",  	 --  2927 	 211 
	 "101110001100",  	 --  2956 	 212 
	 "101110101001",  	 --  2985 	 213 
	 "101111000110",  	 --  3014 	 214 
	 "101111100011",  	 --  3043 	 215 
	 "110000000000",  	 --  3072 	 216 
	 "110000011101",  	 --  3101 	 217 
	 "110000111010",  	 --  3130 	 218 
	 "110001010111",  	 --  3159 	 219 
	 "110001110100",  	 --  3188 	 220 
	 "110010010001",  	 --  3217 	 221 
	 "110010101101",  	 --  3245 	 222 
	 "110011001010",  	 --  3274 	 223 
	 "110011100111",  	 --  3303 	 224 
	 "110100000100",  	 --  3332 	 225 
	 "110100100001",  	 --  3361 	 226 
	 "110100111110",  	 --  3390 	 227 
	 "110101011011",  	 --  3419 	 228 
	 "110101111000",  	 --  3448 	 229 
	 "110110010101",  	 --  3477 	 230 
	 "110110110010",  	 --  3506 	 231 
	 "110111001111",  	 --  3535 	 232 
	 "110111101100",  	 --  3564 	 233 
	 "111000001001",  	 --  3593 	 234 
	 "111000100110",  	 --  3622 	 235 
	 "111001000011",  	 --  3651 	 236 
	 "111001100000",  	 --  3680 	 237 
	 "111001111101",  	 --  3709 	 238 
	 "111010011010",  	 --  3738 	 239 
	 "111010110111",  	 --  3767 	 240 
	 "111011010100",  	 --  3796 	 241 
	 "111011110001",  	 --  3825 	 242 
	 "111100001110",  	 --  3854 	 243 
	 "111100101011",  	 --  3883 	 244 
	 "111101001000",  	 --  3912 	 245 
	 "111101100101",  	 --  3941 	 246 
	 "111110000010",  	 --  3970 	 247 
	 "111110011111",  	 --  3999 	 248 
	 "111110111100",  	 --  4028 	 249 
	 "111111011001",  	 --  4057 	 250 
	 "111111110110",  	 --  4086 	 251 
	 "100011110110",  	 --  2294 	 252 
	 "100100010011",  	 --  2323 	 253 
	 "100100110000",  	 --  2352 	 254 
	 "100101001101",  	 --  2381 	 255 
	 "100101101010",  	 --  2410 	 256 
	 "100110000111",  	 --  2439 	 257 
	 "100110100100",  	 --  2468 	 258 
	 "100111000001",  	 --  2497 	 259 
	 "100111011110",  	 --  2526 	 260 
	 "100111111011",  	 --  2555 	 261 
	 "101000011000",  	 --  2584 	 262 
	 "101000110101",  	 --  2613 	 263 
	 "101001010010",  	 --  2642 	 264 
	 "101001101111",  	 --  2671 	 265 
	 "101010001100",  	 --  2700 	 266 
	 "101010101001",  	 --  2729 	 267 
	 "101011000110",  	 --  2758 	 268 
	 "101011100011",  	 --  2787 	 269 
	 "101100000000",  	 --  2816 	 270 
	 "101100011101",  	 --  2845 	 271 
	 "101100111010",  	 --  2874 	 272 
	 "101101010111",  	 --  2903 	 273 
	 "101101110100",  	 --  2932 	 274 
	 "101110010001",  	 --  2961 	 275 
	 "101110101110",  	 --  2990 	 276 
	 "101111001011",  	 --  3019 	 277 
	 "101111101000",  	 --  3048 	 278 
	 "110000000101",  	 --  3077 	 279 
	 "110000100010",  	 --  3106 	 280 
	 "110000111111",  	 --  3135 	 281 
	 "110001011011",  	 --  3163 	 282 
	 "110001111000",  	 --  3192 	 283 
	 "110010010101",  	 --  3221 	 284 
	 "110010110010",  	 --  3250 	 285 
	 "110011001111",  	 --  3279 	 286 
	 "110011101100",  	 --  3308 	 287 
	 "110100001001",  	 --  3337 	 288 
	 "110100100110",  	 --  3366 	 289 
	 "110101000011",  	 --  3395 	 290 
	 "110101100000",  	 --  3424 	 291 
	 "110101111101",  	 --  3453 	 292 
	 "110110011010",  	 --  3482 	 293 
	 "110110110111",  	 --  3511 	 294 
	 "110111010100",  	 --  3540 	 295 
	 "110111110001",  	 --  3569 	 296 
	 "111000001110",  	 --  3598 	 297 
	 "111000101011",  	 --  3627 	 298 
	 "111001001000",  	 --  3656 	 299 
	 "111001100101",  	 --  3685 	 300 
	 "111010000010",  	 --  3714 	 301 
	 "111010011111",  	 --  3743 	 302 
	 "111010111100",  	 --  3772 	 303 
	 "111011011001",  	 --  3801 	 304 
	 "111011110110",  	 --  3830 	 305 
	 "111100010011",  	 --  3859 	 306 
	 "111100110000",  	 --  3888 	 307 
	 "111101001101",  	 --  3917 	 308 
	 "111101101010",  	 --  3946 	 309 
	 "111110000111",  	 --  3975 	 310 
	 "111110100011",  	 --  4003 	 311 
	 "111111000000",  	 --  4032 	 312 
	 "111111011101",  	 --  4061 	 313 
	 "111111111010",  	 --  4090 	 314 
	 "100011111011",  	 --  2299 	 315 
	 "100100011000",  	 --  2328 	 316 
	 "100100110101",  	 --  2357 	 317 
	 "100101010010",  	 --  2386 	 318 
	 "100101101111",  	 --  2415 	 319 
	 "100110001100",  	 --  2444 	 320 
	 "100110101001",  	 --  2473 	 321 
	 "100111000110",  	 --  2502 	 322 
	 "100111100011",  	 --  2531 	 323 
	 "101000000000",  	 --  2560 	 324 
	 "101000011101",  	 --  2589 	 325 
	 "101000111010",  	 --  2618 	 326 
	 "101001010111",  	 --  2647 	 327 
	 "101001110100",  	 --  2676 	 328 
	 "101010010001",  	 --  2705 	 329 
	 "101010101110",  	 --  2734 	 330 
	 "101011001011",  	 --  2763 	 331 
	 "101011101000",  	 --  2792 	 332 
	 "101100000101",  	 --  2821 	 333 
	 "101100100010",  	 --  2850 	 334 
	 "101100111111",  	 --  2879 	 335 
	 "101101011100",  	 --  2908 	 336 
	 "101101111001",  	 --  2937 	 337 
	 "101110010110",  	 --  2966 	 338 
	 "101110110011",  	 --  2995 	 339 
	 "101111010000",  	 --  3024 	 340 
	 "101111101100",  	 --  3052 	 341 
	 "110000001001",  	 --  3081 	 342 
	 "110000100110",  	 --  3110 	 343 
	 "110001000011",  	 --  3139 	 344 
	 "110001100000",  	 --  3168 	 345 
	 "110001111101",  	 --  3197 	 346 
	 "110010011010",  	 --  3226 	 347 
	 "110010110111",  	 --  3255 	 348 
	 "110011010100",  	 --  3284 	 349 
	 "110011110001",  	 --  3313 	 350 
	 "110100001110",  	 --  3342 	 351 
	 "110100101011",  	 --  3371 	 352 
	 "110101001000",  	 --  3400 	 353 
	 "110101100101",  	 --  3429 	 354 
	 "110110000010",  	 --  3458 	 355 
	 "110110011111",  	 --  3487 	 356 
	 "110110111100",  	 --  3516 	 357 
	 "110111011001",  	 --  3545 	 358 
	 "110111110110",  	 --  3574 	 359 
	 "111000010011",  	 --  3603 	 360 
	 "111000110000",  	 --  3632 	 361 
	 "111001001101",  	 --  3661 	 362 
	 "111001101010",  	 --  3690 	 363 
	 "111010000111",  	 --  3719 	 364 
	 "111010100100",  	 --  3748 	 365 
	 "111011000001",  	 --  3777 	 366 
	 "111011011110",  	 --  3806 	 367 
	 "111011111011",  	 --  3835 	 368 
	 "111100011000",  	 --  3864 	 369 
	 "111100110100",  	 --  3892 	 370 
	 "111101010001",  	 --  3921 	 371 
	 "111101101110",  	 --  3950 	 372 
	 "111110001011",  	 --  3979 	 373 
	 "111110101000",  	 --  4008 	 374 
	 "111111000101",  	 --  4037 	 375 
	 "111111100010",  	 --  4066 	 376 
	 "100011100011",  	 --  2275 	 377 
	 "100100000000",  	 --  2304 	 378 
	 "100100011101",  	 --  2333 	 379 
	 "100100111010",  	 --  2362 	 380 
	 "100101010111",  	 --  2391 	 381 
	 "100101110100",  	 --  2420 	 382 
	 "100110010001",  	 --  2449 	 383 
	 "100110101110",  	 --  2478 	 384 
	 "100111001011",  	 --  2507 	 385 
	 "100111101000",  	 --  2536 	 386 
	 "101000000101",  	 --  2565 	 387 
	 "101000100010",  	 --  2594 	 388 
	 "101000111111",  	 --  2623 	 389 
	 "101001011100",  	 --  2652 	 390 
	 "101001111001",  	 --  2681 	 391 
	 "101010010110",  	 --  2710 	 392 
	 "101010110011",  	 --  2739 	 393 
	 "101011010000",  	 --  2768 	 394 
	 "101011101101",  	 --  2797 	 395 
	 "101100001010",  	 --  2826 	 396 
	 "101100100111",  	 --  2855 	 397 
	 "101101000100",  	 --  2884 	 398 
	 "101101100001",  	 --  2913 	 399 
	 "101101111101",  	 --  2941 	 400 
	 "101110011010",  	 --  2970 	 401 
	 "101110110111",  	 --  2999 	 402 
	 "101111010100",  	 --  3028 	 403 
	 "101111110001",  	 --  3057 	 404 
	 "110000001110",  	 --  3086 	 405 
	 "110000101011",  	 --  3115 	 406 
	 "110001001000",  	 --  3144 	 407 
	 "110001100101",  	 --  3173 	 408 
	 "110010000010",  	 --  3202 	 409 
	 "110010011111",  	 --  3231 	 410 
	 "110010111100",  	 --  3260 	 411 
	 "110011011001",  	 --  3289 	 412 
	 "110011110110",  	 --  3318 	 413 
	 "110100010011",  	 --  3347 	 414 
	 "110100110000",  	 --  3376 	 415 
	 "110101001101",  	 --  3405 	 416 
	 "110101101010",  	 --  3434 	 417 
	 "110110000111",  	 --  3463 	 418 
	 "110110100100",  	 --  3492 	 419 
	 "110111000001",  	 --  3521 	 420 
	 "110111011110",  	 --  3550 	 421 
	 "110111111011",  	 --  3579 	 422 
	 "111000011000",  	 --  3608 	 423 
	 "111000110101",  	 --  3637 	 424 
	 "111001010010",  	 --  3666 	 425 
	 "111001101111",  	 --  3695 	 426 
	 "111010001100",  	 --  3724 	 427 
	 "111010101001",  	 --  3753 	 428 
	 "111011000101",  	 --  3781 	 429 
	 "111011100010",  	 --  3810 	 430 
	 "111011111111",  	 --  3839 	 431 
	 "111100011100",  	 --  3868 	 432 
	 "111100111001",  	 --  3897 	 433 
	 "111101010110",  	 --  3926 	 434 
	 "111101110011",  	 --  3955 	 435 
	 "111110010000",  	 --  3984 	 436 
	 "111110101101",  	 --  4013 	 437 
	 "111111001010",  	 --  4042 	 438 
	 "111111100111",  	 --  4071 	 439 
	 "100011101000",  	 --  2280 	 440 
	 "100100000101",  	 --  2309 	 441 
	 "100100100010",  	 --  2338 	 442 
	 "100100111111",  	 --  2367 	 443 
	 "100101011100",  	 --  2396 	 444 
	 "100101111001",  	 --  2425 	 445 
	 "100110010110",  	 --  2454 	 446 
	 "100110110011",  	 --  2483 	 447 
	 "100111010000",  	 --  2512 	 448 
	 "100111101101",  	 --  2541 	 449 
	 "101000001010",  	 --  2570 	 450 
	 "101000100111",  	 --  2599 	 451 
	 "101001000100",  	 --  2628 	 452 
	 "101001100001",  	 --  2657 	 453 
	 "101001111110",  	 --  2686 	 454 
	 "101010011011",  	 --  2715 	 455 
	 "101010111000",  	 --  2744 	 456 
	 "101011010101",  	 --  2773 	 457 
	 "101011110010",  	 --  2802 	 458 
	 "101100001110",  	 --  2830 	 459 
	 "101100101011",  	 --  2859 	 460 
	 "101101001000",  	 --  2888 	 461 
	 "101101100101",  	 --  2917 	 462 
	 "101110000010",  	 --  2946 	 463 
	 "101110011111",  	 --  2975 	 464 
	 "101110111100",  	 --  3004 	 465 
	 "101111011001",  	 --  3033 	 466 
	 "101111110110",  	 --  3062 	 467 
	 "110000010011",  	 --  3091 	 468 
	 "110000110000",  	 --  3120 	 469 
	 "110001001101",  	 --  3149 	 470 
	 "110001101010",  	 --  3178 	 471 
	 "110010000111",  	 --  3207 	 472 
	 "110010100100",  	 --  3236 	 473 
	 "110011000001",  	 --  3265 	 474 
	 "110011011110",  	 --  3294 	 475 
	 "110011111011",  	 --  3323 	 476 
	 "110100011000",  	 --  3352 	 477 
	 "110100110101",  	 --  3381 	 478 
	 "110101010010",  	 --  3410 	 479 
	 "110101101111",  	 --  3439 	 480 
	 "110110001100",  	 --  3468 	 481 
	 "110110101001",  	 --  3497 	 482 
	 "110111000110",  	 --  3526 	 483 
	 "110111100011",  	 --  3555 	 484 
	 "111000000000",  	 --  3584 	 485 
	 "111000011101",  	 --  3613 	 486 
	 "111000111010",  	 --  3642 	 487 
	 "111001010111",  	 --  3671 	 488 
	 "111001110011",  	 --  3699 	 489 
	 "111010010000",  	 --  3728 	 490 
	 "111010101101",  	 --  3757 	 491 
	 "111011001010",  	 --  3786 	 492 
	 "111011100111",  	 --  3815 	 493 
	 "111100000100",  	 --  3844 	 494 
	 "111100100001",  	 --  3873 	 495 
	 "111100111110",  	 --  3902 	 496 
	 "111101011011",  	 --  3931 	 497 
	 "111101111000",  	 --  3960 	 498 
	 "111110010101",  	 --  3989 	 499 
	 "111110110010",  	 --  4018 	 500 
	 "111111001111",  	 --  4047 	 501 
	 "111111101100",  	 --  4076 	 502 
	 "100011101101",  	 --  2285 	 503 
	 "100100001010",  	 --  2314 	 504 
	 "100100100111",  	 --  2343 	 505 
	 "100101000100",  	 --  2372 	 506 
	 "100101100001",  	 --  2401 	 507 
	 "100101111110",  	 --  2430 	 508 
	 "100110011011",  	 --  2459 	 509 
	 "100110111000",  	 --  2488 	 510 
 	"100111010101");  --  2517 	 511
	begin 
		return tmp;
	end init_rom;
	signal rom : memory_t := init_rom;
begin
	process(clk,ADDR)
		variable addr2 : natural range 0 to 2**m - 1;
	begin
	addr2 := to_integer(unsigned(ADDR));
	if( falling_edge(clk)) then
		q <= rom(addr2);
	end if;
	end process;
end rtl;
