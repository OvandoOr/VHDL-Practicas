library IEEE;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;

entity Comparador_MenorIgual is
	generic(
	n: integer := 8
	);
	port(
	A: 		in std_logic_vector(n-1 downto 0);
	B:		in std_logic_vector(n-1 downto 0);
	MenorIgual:	out std_logic
	);
end Comparador_MenorIgual;

architecture Comparador of Comparador_MenorIgual is
begin
	combinacional: process(A,B)
	begin
		if(A <= B) then
			MenorIgual <= '1';
		else
			MenorIgual <= '0';
		end if;
	end process combinacional;

end Comparador;


















































































































































































































































































































































































































































































































































































